magic
tech sky130A
magscale 1 2
timestamp 1763265783
<< obsli1 >>
rect 1104 2159 9292 10353
<< obsm1 >>
rect 14 2128 10382 10384
<< metal2 >>
rect 1306 11817 1362 12617
rect 3882 11817 3938 12617
rect 6458 11817 6514 12617
rect 9034 11817 9090 12617
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 7746 0 7802 800
rect 10322 0 10378 800
<< obsm2 >>
rect 20 11761 1250 11817
rect 1418 11761 3826 11817
rect 3994 11761 6402 11817
rect 6570 11761 8978 11817
rect 9146 11761 10376 11817
rect 20 856 10376 11761
rect 130 800 2538 856
rect 2706 800 5114 856
rect 5282 800 7690 856
rect 7858 800 10266 856
<< metal3 >>
rect 0 10888 800 11008
rect 9673 10888 10473 11008
rect 0 8168 800 8288
rect 9673 8168 10473 8288
rect 0 5448 800 5568
rect 9673 5448 10473 5568
rect 0 2728 800 2848
rect 9673 2728 10473 2848
<< obsm3 >>
rect 880 10808 9593 10981
rect 800 8368 9673 10808
rect 880 8088 9593 8368
rect 800 5648 9673 8088
rect 880 5368 9593 5648
rect 800 2928 9673 5368
rect 880 2648 9593 2928
rect 800 2143 9673 2648
<< metal4 >>
rect 1967 2128 2287 10384
rect 2627 2128 2947 10384
rect 4014 2128 4334 10384
rect 4674 2128 4994 10384
rect 6061 2128 6381 10384
rect 6721 2128 7041 10384
rect 8108 2128 8428 10384
rect 8768 2128 9088 10384
<< metal5 >>
rect 1056 9816 9340 10136
rect 1056 9156 9340 9476
rect 1056 7776 9340 8096
rect 1056 7116 9340 7436
rect 1056 5736 9340 6056
rect 1056 5076 9340 5396
rect 1056 3696 9340 4016
rect 1056 3036 9340 3356
<< labels >>
rlabel metal3 s 9673 8168 10473 8288 6 A[0]
port 1 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 A[2]
port 3 nsew signal input
rlabel metal2 s 6458 11817 6514 12617 6 A[3]
port 4 nsew signal input
rlabel metal2 s 3882 11817 3938 12617 6 B[0]
port 5 nsew signal input
rlabel metal2 s 18 0 74 800 6 B[1]
port 6 nsew signal input
rlabel metal3 s 9673 10888 10473 11008 6 B[2]
port 7 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 B[3]
port 8 nsew signal input
rlabel metal4 s 2627 2128 2947 10384 6 VGND
port 9 nsew ground bidirectional
rlabel metal4 s 4674 2128 4994 10384 6 VGND
port 9 nsew ground bidirectional
rlabel metal4 s 6721 2128 7041 10384 6 VGND
port 9 nsew ground bidirectional
rlabel metal4 s 8768 2128 9088 10384 6 VGND
port 9 nsew ground bidirectional
rlabel metal5 s 1056 3696 9340 4016 6 VGND
port 9 nsew ground bidirectional
rlabel metal5 s 1056 5736 9340 6056 6 VGND
port 9 nsew ground bidirectional
rlabel metal5 s 1056 7776 9340 8096 6 VGND
port 9 nsew ground bidirectional
rlabel metal5 s 1056 9816 9340 10136 6 VGND
port 9 nsew ground bidirectional
rlabel metal4 s 1967 2128 2287 10384 6 VPWR
port 10 nsew power bidirectional
rlabel metal4 s 4014 2128 4334 10384 6 VPWR
port 10 nsew power bidirectional
rlabel metal4 s 6061 2128 6381 10384 6 VPWR
port 10 nsew power bidirectional
rlabel metal4 s 8108 2128 8428 10384 6 VPWR
port 10 nsew power bidirectional
rlabel metal5 s 1056 3036 9340 3356 6 VPWR
port 10 nsew power bidirectional
rlabel metal5 s 1056 5076 9340 5396 6 VPWR
port 10 nsew power bidirectional
rlabel metal5 s 1056 7116 9340 7436 6 VPWR
port 10 nsew power bidirectional
rlabel metal5 s 1056 9156 9340 9476 6 VPWR
port 10 nsew power bidirectional
rlabel metal2 s 2594 0 2650 800 6 clk
port 11 nsew signal input
rlabel metal3 s 9673 2728 10473 2848 6 result[0]
port 12 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 result[1]
port 13 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 result[2]
port 14 nsew signal output
rlabel metal2 s 9034 11817 9090 12617 6 result[3]
port 15 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 rst
port 16 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 sel[0]
port 17 nsew signal input
rlabel metal2 s 1306 11817 1362 12617 6 sel[1]
port 18 nsew signal input
rlabel metal3 s 9673 5448 10473 5568 6 sel[2]
port 19 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10473 12617
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 517278
string GDS_FILE /openlane/designs/alu4bit/runs/RUN_2025.11.16_04.02.04/results/signoff/alu4bit.magic.gds
string GDS_START 251122
<< end >>

