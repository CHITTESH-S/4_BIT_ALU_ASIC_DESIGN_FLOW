magic
tech sky130A
magscale 1 2
timestamp 1763265782
<< viali >>
rect 8217 10217 8251 10251
rect 1593 10149 1627 10183
rect 1409 10013 1443 10047
rect 1777 10013 1811 10047
rect 4077 10013 4111 10047
rect 6653 10013 6687 10047
rect 8677 10013 8711 10047
rect 4261 9945 4295 9979
rect 8309 9945 8343 9979
rect 1961 9877 1995 9911
rect 6745 9877 6779 9911
rect 8585 9877 8619 9911
rect 4905 9673 4939 9707
rect 3341 9605 3375 9639
rect 6101 9605 6135 9639
rect 8553 9605 8587 9639
rect 8769 9605 8803 9639
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 2973 9537 3007 9571
rect 3249 9537 3283 9571
rect 3525 9537 3559 9571
rect 3801 9537 3835 9571
rect 4077 9537 4111 9571
rect 4629 9537 4663 9571
rect 4721 9537 4755 9571
rect 5641 9537 5675 9571
rect 5825 9537 5859 9571
rect 6009 9537 6043 9571
rect 6193 9547 6227 9581
rect 6561 9537 6595 9571
rect 6745 9537 6779 9571
rect 7205 9537 7239 9571
rect 7389 9537 7423 9571
rect 7481 9537 7515 9571
rect 8125 9537 8159 9571
rect 8309 9537 8343 9571
rect 3157 9469 3191 9503
rect 4353 9469 4387 9503
rect 4905 9469 4939 9503
rect 7021 9469 7055 9503
rect 7757 9469 7791 9503
rect 3249 9401 3283 9435
rect 4261 9401 4295 9435
rect 6377 9401 6411 9435
rect 7849 9401 7883 9435
rect 2881 9333 2915 9367
rect 3709 9333 3743 9367
rect 4169 9333 4203 9367
rect 5733 9333 5767 9367
rect 8401 9333 8435 9367
rect 8585 9333 8619 9367
rect 7757 9129 7791 9163
rect 2881 8993 2915 9027
rect 2789 8925 2823 8959
rect 4721 8925 4755 8959
rect 4905 8925 4939 8959
rect 4997 8925 5031 8959
rect 5089 8925 5123 8959
rect 5641 8925 5675 8959
rect 5825 8925 5859 8959
rect 6009 8925 6043 8959
rect 6101 8925 6135 8959
rect 7573 8925 7607 8959
rect 5365 8857 5399 8891
rect 5733 8857 5767 8891
rect 7389 8857 7423 8891
rect 3157 8789 3191 8823
rect 5457 8789 5491 8823
rect 8953 8585 8987 8619
rect 1409 8449 1443 8483
rect 7829 8449 7863 8483
rect 7573 8381 7607 8415
rect 1593 8245 1627 8279
rect 3341 8041 3375 8075
rect 3801 8041 3835 8075
rect 5549 8041 5583 8075
rect 5641 8041 5675 8075
rect 3433 7973 3467 8007
rect 2789 7905 2823 7939
rect 2973 7837 3007 7871
rect 3433 7837 3467 7871
rect 4077 7837 4111 7871
rect 5181 7837 5215 7871
rect 5641 7837 5675 7871
rect 8677 7837 8711 7871
rect 2544 7769 2578 7803
rect 3801 7769 3835 7803
rect 3985 7769 4019 7803
rect 8493 7769 8527 7803
rect 1409 7701 1443 7735
rect 3065 7701 3099 7735
rect 3157 7701 3191 7735
rect 5273 7701 5307 7735
rect 5365 7701 5399 7735
rect 2513 7497 2547 7531
rect 3065 7497 3099 7531
rect 5365 7497 5399 7531
rect 6377 7497 6411 7531
rect 7665 7429 7699 7463
rect 7881 7429 7915 7463
rect 2053 7361 2087 7395
rect 2145 7361 2179 7395
rect 2237 7361 2271 7395
rect 2329 7361 2363 7395
rect 4353 7361 4387 7395
rect 5549 7361 5583 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 5917 7361 5951 7395
rect 6745 7361 6779 7395
rect 6653 7293 6687 7327
rect 7849 7157 7883 7191
rect 8033 7157 8067 7191
rect 3249 6953 3283 6987
rect 5549 6953 5583 6987
rect 8125 6953 8159 6987
rect 4470 6817 4504 6851
rect 7389 6817 7423 6851
rect 7481 6817 7515 6851
rect 2973 6749 3007 6783
rect 3985 6749 4019 6783
rect 5733 6749 5767 6783
rect 5825 6749 5859 6783
rect 7021 6749 7055 6783
rect 7159 6749 7193 6783
rect 7849 6749 7883 6783
rect 7941 6749 7975 6783
rect 8217 6749 8251 6783
rect 8309 6749 8343 6783
rect 8493 6749 8527 6783
rect 3249 6681 3283 6715
rect 4353 6681 4387 6715
rect 5549 6681 5583 6715
rect 3065 6613 3099 6647
rect 4261 6613 4295 6647
rect 4629 6613 4663 6647
rect 7021 6613 7055 6647
rect 8677 6613 8711 6647
rect 1777 6409 1811 6443
rect 2815 6409 2849 6443
rect 3709 6409 3743 6443
rect 4813 6409 4847 6443
rect 8033 6409 8067 6443
rect 2053 6341 2087 6375
rect 2605 6341 2639 6375
rect 3985 6341 4019 6375
rect 5181 6341 5215 6375
rect 1961 6273 1995 6307
rect 3888 6273 3922 6307
rect 4077 6273 4111 6307
rect 4260 6273 4294 6307
rect 4353 6273 4387 6307
rect 4721 6273 4755 6307
rect 4997 6273 5031 6307
rect 5457 6273 5491 6307
rect 5733 6273 5767 6307
rect 7665 6273 7699 6307
rect 7757 6273 7791 6307
rect 7849 6273 7883 6307
rect 8585 6273 8619 6307
rect 2513 6205 2547 6239
rect 5089 6205 5123 6239
rect 5273 6205 5307 6239
rect 2329 6137 2363 6171
rect 2973 6137 3007 6171
rect 8125 6137 8159 6171
rect 2789 6069 2823 6103
rect 5641 6069 5675 6103
rect 8309 6069 8343 6103
rect 4353 5865 4387 5899
rect 4445 5797 4479 5831
rect 4997 5797 5031 5831
rect 6561 5797 6595 5831
rect 7849 5797 7883 5831
rect 3893 5729 3927 5763
rect 1501 5661 1535 5695
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 4169 5661 4203 5695
rect 4435 5661 4469 5695
rect 4721 5661 4755 5695
rect 5181 5661 5215 5695
rect 7205 5661 7239 5695
rect 7297 5661 7331 5695
rect 7481 5661 7515 5695
rect 8769 5661 8803 5695
rect 5273 5593 5307 5627
rect 1593 5525 1627 5559
rect 4629 5525 4663 5559
rect 8585 5525 8619 5559
rect 2237 5321 2271 5355
rect 2697 5321 2731 5355
rect 3617 5321 3651 5355
rect 5641 5321 5675 5355
rect 7573 5321 7607 5355
rect 3433 5253 3467 5287
rect 5181 5253 5215 5287
rect 5273 5253 5307 5287
rect 1869 5185 1903 5219
rect 2876 5185 2910 5219
rect 2973 5185 3007 5219
rect 3065 5185 3099 5219
rect 3248 5185 3282 5219
rect 3341 5185 3375 5219
rect 3709 5185 3743 5219
rect 4997 5185 5031 5219
rect 5365 5185 5399 5219
rect 5917 5185 5951 5219
rect 6193 5185 6227 5219
rect 7941 5185 7975 5219
rect 8677 5185 8711 5219
rect 7849 5117 7883 5151
rect 8217 5117 8251 5151
rect 2421 5049 2455 5083
rect 2237 4981 2271 5015
rect 3433 4981 3467 5015
rect 5549 4981 5583 5015
rect 5825 4981 5859 5015
rect 8493 4981 8527 5015
rect 3801 4777 3835 4811
rect 5825 4777 5859 4811
rect 6193 4777 6227 4811
rect 4445 4709 4479 4743
rect 4261 4641 4295 4675
rect 3985 4573 4019 4607
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 5733 4573 5767 4607
rect 4629 4437 4663 4471
rect 5733 4165 5767 4199
rect 5917 4165 5951 4199
rect 6009 4097 6043 4131
rect 6137 4097 6171 4131
rect 6562 4097 6596 4131
rect 6653 4097 6687 4131
rect 6929 4097 6963 4131
rect 5917 4029 5951 4063
rect 6837 4029 6871 4063
rect 6377 3893 6411 3927
rect 2421 3689 2455 3723
rect 3249 3689 3283 3723
rect 5641 3689 5675 3723
rect 5825 3553 5859 3587
rect 2421 3485 2455 3519
rect 2605 3485 2639 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4169 3485 4203 3519
rect 4279 3485 4313 3519
rect 4445 3485 4479 3519
rect 4813 3485 4847 3519
rect 5273 3485 5307 3519
rect 5549 3485 5583 3519
rect 1501 3417 1535 3451
rect 3157 3417 3191 3451
rect 1593 3349 1627 3383
rect 2789 3349 2823 3383
rect 3801 3349 3835 3383
rect 5181 3349 5215 3383
rect 6101 3349 6135 3383
rect 1593 3145 1627 3179
rect 4629 3145 4663 3179
rect 6745 3145 6779 3179
rect 7113 3145 7147 3179
rect 8585 3145 8619 3179
rect 4353 3077 4387 3111
rect 5917 3077 5951 3111
rect 6377 3077 6411 3111
rect 7450 3077 7484 3111
rect 1501 3009 1535 3043
rect 4445 3009 4479 3043
rect 4721 3009 4755 3043
rect 5549 3009 5583 3043
rect 6561 3009 6595 3043
rect 6837 3009 6871 3043
rect 6929 2993 6963 3027
rect 7205 3009 7239 3043
rect 8677 3009 8711 3043
rect 3065 2873 3099 2907
rect 6101 2873 6135 2907
rect 4445 2805 4479 2839
rect 5917 2805 5951 2839
rect 8861 2805 8895 2839
rect 1409 2601 1443 2635
rect 4169 2601 4203 2635
rect 5457 2601 5491 2635
rect 7849 2601 7883 2635
rect 8585 2601 8619 2635
rect 2789 2465 2823 2499
rect 3801 2397 3835 2431
rect 3893 2397 3927 2431
rect 4261 2397 4295 2431
rect 5273 2397 5307 2431
rect 8033 2397 8067 2431
rect 8769 2397 8803 2431
rect 2544 2329 2578 2363
rect 3985 2261 4019 2295
rect 4261 2261 4295 2295
<< metal1 >>
rect 1104 10362 9292 10384
rect 1104 10310 1973 10362
rect 2025 10310 2037 10362
rect 2089 10310 2101 10362
rect 2153 10310 2165 10362
rect 2217 10310 2229 10362
rect 2281 10310 4020 10362
rect 4072 10310 4084 10362
rect 4136 10310 4148 10362
rect 4200 10310 4212 10362
rect 4264 10310 4276 10362
rect 4328 10310 6067 10362
rect 6119 10310 6131 10362
rect 6183 10310 6195 10362
rect 6247 10310 6259 10362
rect 6311 10310 6323 10362
rect 6375 10310 8114 10362
rect 8166 10310 8178 10362
rect 8230 10310 8242 10362
rect 8294 10310 8306 10362
rect 8358 10310 8370 10362
rect 8422 10310 9292 10362
rect 1104 10288 9292 10310
rect 1302 10208 1308 10260
rect 1360 10208 1366 10260
rect 8205 10251 8263 10257
rect 8205 10217 8217 10251
rect 8251 10248 8263 10251
rect 9030 10248 9036 10260
rect 8251 10220 9036 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 1320 10112 1348 10208
rect 1581 10183 1639 10189
rect 1581 10149 1593 10183
rect 1627 10180 1639 10183
rect 2958 10180 2964 10192
rect 1627 10152 2964 10180
rect 1627 10149 1639 10152
rect 1581 10143 1639 10149
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 1320 10084 1808 10112
rect 934 10004 940 10056
rect 992 10044 998 10056
rect 1780 10053 1808 10084
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 992 10016 1409 10044
rect 992 10004 998 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 3936 10016 4077 10044
rect 3936 10004 3942 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6641 10047 6699 10053
rect 6641 10044 6653 10047
rect 6512 10016 6653 10044
rect 6512 10004 6518 10016
rect 6641 10013 6653 10016
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10044 8723 10047
rect 9214 10044 9220 10056
rect 8711 10016 9220 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 4249 9979 4307 9985
rect 4249 9945 4261 9979
rect 4295 9976 4307 9979
rect 7098 9976 7104 9988
rect 4295 9948 7104 9976
rect 4295 9945 4307 9948
rect 4249 9939 4307 9945
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 8297 9979 8355 9985
rect 8297 9945 8309 9979
rect 8343 9976 8355 9979
rect 8478 9976 8484 9988
rect 8343 9948 8484 9976
rect 8343 9945 8355 9948
rect 8297 9939 8355 9945
rect 8478 9936 8484 9948
rect 8536 9936 8542 9988
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 1949 9911 2007 9917
rect 1949 9908 1961 9911
rect 1912 9880 1961 9908
rect 1912 9868 1918 9880
rect 1949 9877 1961 9880
rect 1995 9877 2007 9911
rect 1949 9871 2007 9877
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6696 9880 6745 9908
rect 6696 9868 6702 9880
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 1104 9818 9292 9840
rect 1104 9766 2633 9818
rect 2685 9766 2697 9818
rect 2749 9766 2761 9818
rect 2813 9766 2825 9818
rect 2877 9766 2889 9818
rect 2941 9766 4680 9818
rect 4732 9766 4744 9818
rect 4796 9766 4808 9818
rect 4860 9766 4872 9818
rect 4924 9766 4936 9818
rect 4988 9766 6727 9818
rect 6779 9766 6791 9818
rect 6843 9766 6855 9818
rect 6907 9766 6919 9818
rect 6971 9766 6983 9818
rect 7035 9766 8774 9818
rect 8826 9766 8838 9818
rect 8890 9766 8902 9818
rect 8954 9766 8966 9818
rect 9018 9766 9030 9818
rect 9082 9766 9292 9818
rect 1104 9744 9292 9766
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3016 9676 3556 9704
rect 3016 9664 3022 9676
rect 3329 9639 3387 9645
rect 3329 9636 3341 9639
rect 2700 9608 3341 9636
rect 2700 9577 2728 9608
rect 3329 9605 3341 9608
rect 3375 9605 3387 9639
rect 3329 9599 3387 9605
rect 3528 9636 3556 9676
rect 4890 9664 4896 9716
rect 4948 9664 4954 9716
rect 5552 9676 6316 9704
rect 3878 9636 3884 9648
rect 3528 9608 3884 9636
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 2884 9500 2912 9531
rect 2958 9528 2964 9580
rect 3016 9528 3022 9580
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3418 9568 3424 9580
rect 3283 9540 3424 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 3528 9577 3556 9608
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 5552 9636 5580 9676
rect 6089 9639 6147 9645
rect 6089 9636 6101 9639
rect 4080 9608 5580 9636
rect 5644 9608 6101 9636
rect 4080 9577 4108 9608
rect 5644 9580 5672 9608
rect 6089 9605 6101 9608
rect 6135 9605 6147 9639
rect 6288 9636 6316 9676
rect 7742 9636 7748 9648
rect 6288 9608 7144 9636
rect 6089 9599 6147 9605
rect 6181 9581 6239 9587
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3835 9540 4077 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 3145 9503 3203 9509
rect 2884 9472 3004 9500
rect 2866 9324 2872 9376
rect 2924 9324 2930 9376
rect 2976 9364 3004 9472
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3804 9500 3832 9531
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4212 9540 4476 9568
rect 4212 9528 4218 9540
rect 3191 9472 3832 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 4341 9503 4399 9509
rect 4341 9500 4353 9503
rect 3936 9472 4353 9500
rect 3936 9460 3942 9472
rect 4341 9469 4353 9472
rect 4387 9469 4399 9503
rect 4448 9500 4476 9540
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 4617 9571 4675 9577
rect 4617 9568 4629 9571
rect 4580 9540 4629 9568
rect 4580 9528 4586 9540
rect 4617 9537 4629 9540
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4755 9540 5028 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4724 9500 4752 9531
rect 4448 9472 4752 9500
rect 4893 9503 4951 9509
rect 4341 9463 4399 9469
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 3237 9435 3295 9441
rect 3237 9401 3249 9435
rect 3283 9432 3295 9435
rect 4062 9432 4068 9444
rect 3283 9404 4068 9432
rect 3283 9401 3295 9404
rect 3237 9395 3295 9401
rect 3252 9364 3280 9395
rect 4062 9392 4068 9404
rect 4120 9392 4126 9444
rect 4249 9435 4307 9441
rect 4249 9401 4261 9435
rect 4295 9432 4307 9435
rect 4614 9432 4620 9444
rect 4295 9404 4620 9432
rect 4295 9401 4307 9404
rect 4249 9395 4307 9401
rect 4614 9392 4620 9404
rect 4672 9432 4678 9444
rect 4908 9432 4936 9463
rect 5000 9444 5028 9540
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 5859 9540 5948 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 5920 9444 5948 9540
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6181 9547 6193 9581
rect 6227 9578 6239 9581
rect 6227 9550 6316 9578
rect 6227 9547 6239 9550
rect 6181 9541 6239 9547
rect 6288 9500 6316 9550
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6420 9540 6561 9568
rect 6420 9528 6426 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6748 9500 6776 9531
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6288 9472 7021 9500
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 4672 9404 4936 9432
rect 4672 9392 4678 9404
rect 4982 9392 4988 9444
rect 5040 9392 5046 9444
rect 5092 9404 5856 9432
rect 2976 9336 3280 9364
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3476 9336 3709 9364
rect 3476 9324 3482 9336
rect 3697 9333 3709 9336
rect 3743 9364 3755 9367
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 3743 9336 4169 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 4157 9333 4169 9336
rect 4203 9364 4215 9367
rect 5092 9364 5120 9404
rect 4203 9336 5120 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 5718 9324 5724 9376
rect 5776 9324 5782 9376
rect 5828 9364 5856 9404
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 6365 9435 6423 9441
rect 6365 9432 6377 9435
rect 5960 9404 6377 9432
rect 5960 9392 5966 9404
rect 6365 9401 6377 9404
rect 6411 9401 6423 9435
rect 7116 9432 7144 9608
rect 7392 9608 7748 9636
rect 7392 9577 7420 9608
rect 7742 9596 7748 9608
rect 7800 9636 7806 9648
rect 8541 9639 8599 9645
rect 8541 9636 8553 9639
rect 7800 9608 8553 9636
rect 7800 9596 7806 9608
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7208 9500 7236 9531
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7524 9540 7788 9568
rect 7524 9528 7530 9540
rect 7650 9500 7656 9512
rect 7208 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 7760 9509 7788 9540
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8312 9577 8340 9608
rect 8541 9605 8553 9608
rect 8587 9605 8599 9639
rect 8541 9599 8599 9605
rect 8757 9639 8815 9645
rect 8757 9605 8769 9639
rect 8803 9605 8815 9639
rect 8757 9599 8815 9605
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7892 9540 8125 9568
rect 7892 9528 7898 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 7116 9404 7849 9432
rect 6365 9395 6423 9401
rect 7837 9401 7849 9404
rect 7883 9401 7895 9435
rect 8128 9432 8156 9531
rect 8570 9460 8576 9512
rect 8628 9500 8634 9512
rect 8772 9500 8800 9599
rect 8628 9472 8800 9500
rect 8628 9460 8634 9472
rect 8128 9404 8616 9432
rect 7837 9395 7895 9401
rect 8588 9373 8616 9404
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 5828 9336 8401 9364
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8389 9327 8447 9333
rect 8573 9367 8631 9373
rect 8573 9333 8585 9367
rect 8619 9333 8631 9367
rect 8573 9327 8631 9333
rect 1104 9274 9292 9296
rect 1104 9222 1973 9274
rect 2025 9222 2037 9274
rect 2089 9222 2101 9274
rect 2153 9222 2165 9274
rect 2217 9222 2229 9274
rect 2281 9222 4020 9274
rect 4072 9222 4084 9274
rect 4136 9222 4148 9274
rect 4200 9222 4212 9274
rect 4264 9222 4276 9274
rect 4328 9222 6067 9274
rect 6119 9222 6131 9274
rect 6183 9222 6195 9274
rect 6247 9222 6259 9274
rect 6311 9222 6323 9274
rect 6375 9222 8114 9274
rect 8166 9222 8178 9274
rect 8230 9222 8242 9274
rect 8294 9222 8306 9274
rect 8358 9222 8370 9274
rect 8422 9222 9292 9274
rect 1104 9200 9292 9222
rect 2866 9120 2872 9172
rect 2924 9120 2930 9172
rect 4614 9120 4620 9172
rect 4672 9120 4678 9172
rect 4890 9120 4896 9172
rect 4948 9120 4954 9172
rect 5902 9120 5908 9172
rect 5960 9120 5966 9172
rect 7742 9120 7748 9172
rect 7800 9120 7806 9172
rect 2884 9033 2912 9120
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8956 2835 8959
rect 4632 8956 4660 9120
rect 4908 9092 4936 9120
rect 4908 9064 5856 9092
rect 5718 9024 5724 9036
rect 4908 8996 5724 9024
rect 4908 8965 4936 8996
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 2823 8928 4568 8956
rect 4632 8928 4721 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 4540 8900 4568 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 4982 8916 4988 8968
rect 5040 8916 5046 8968
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5123 8928 5212 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 4522 8848 4528 8900
rect 4580 8888 4586 8900
rect 5184 8888 5212 8928
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 5828 8965 5856 9064
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 4580 8860 5212 8888
rect 4580 8848 4586 8860
rect 5184 8832 5212 8860
rect 5353 8891 5411 8897
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 5721 8891 5779 8897
rect 5399 8860 5672 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 3142 8780 3148 8832
rect 3200 8780 3206 8832
rect 5166 8780 5172 8832
rect 5224 8780 5230 8832
rect 5442 8780 5448 8832
rect 5500 8780 5506 8832
rect 5644 8820 5672 8860
rect 5721 8857 5733 8891
rect 5767 8888 5779 8891
rect 5920 8888 5948 9120
rect 7466 9052 7472 9104
rect 7524 9092 7530 9104
rect 8570 9092 8576 9104
rect 7524 9064 8576 9092
rect 7524 9052 7530 9064
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6454 8956 6460 8968
rect 6135 8928 6460 8956
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 5767 8860 5948 8888
rect 5767 8857 5779 8860
rect 5721 8851 5779 8857
rect 6012 8820 6040 8919
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7282 8956 7288 8968
rect 7156 8928 7288 8956
rect 7156 8916 7162 8928
rect 7282 8916 7288 8928
rect 7340 8956 7346 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7340 8928 7573 8956
rect 7340 8916 7346 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7374 8848 7380 8900
rect 7432 8848 7438 8900
rect 5644 8792 6040 8820
rect 1104 8730 9292 8752
rect 1104 8678 2633 8730
rect 2685 8678 2697 8730
rect 2749 8678 2761 8730
rect 2813 8678 2825 8730
rect 2877 8678 2889 8730
rect 2941 8678 4680 8730
rect 4732 8678 4744 8730
rect 4796 8678 4808 8730
rect 4860 8678 4872 8730
rect 4924 8678 4936 8730
rect 4988 8678 6727 8730
rect 6779 8678 6791 8730
rect 6843 8678 6855 8730
rect 6907 8678 6919 8730
rect 6971 8678 6983 8730
rect 7035 8678 8774 8730
rect 8826 8678 8838 8730
rect 8890 8678 8902 8730
rect 8954 8678 8966 8730
rect 9018 8678 9030 8730
rect 9082 8678 9292 8730
rect 1104 8656 9292 8678
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8536 8588 8953 8616
rect 8536 8576 8542 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 5166 8508 5172 8560
rect 5224 8548 5230 8560
rect 7098 8548 7104 8560
rect 5224 8520 7104 8548
rect 5224 8508 5230 8520
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7817 8483 7875 8489
rect 7817 8480 7829 8483
rect 6972 8452 7829 8480
rect 6972 8440 6978 8452
rect 7817 8449 7829 8452
rect 7863 8449 7875 8483
rect 7817 8443 7875 8449
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 7561 8375 7619 8381
rect 1578 8236 1584 8288
rect 1636 8236 1642 8288
rect 3234 8236 3240 8288
rect 3292 8276 3298 8288
rect 7576 8276 7604 8375
rect 3292 8248 7604 8276
rect 3292 8236 3298 8248
rect 1104 8186 9292 8208
rect 1104 8134 1973 8186
rect 2025 8134 2037 8186
rect 2089 8134 2101 8186
rect 2153 8134 2165 8186
rect 2217 8134 2229 8186
rect 2281 8134 4020 8186
rect 4072 8134 4084 8186
rect 4136 8134 4148 8186
rect 4200 8134 4212 8186
rect 4264 8134 4276 8186
rect 4328 8134 6067 8186
rect 6119 8134 6131 8186
rect 6183 8134 6195 8186
rect 6247 8134 6259 8186
rect 6311 8134 6323 8186
rect 6375 8134 8114 8186
rect 8166 8134 8178 8186
rect 8230 8134 8242 8186
rect 8294 8134 8306 8186
rect 8358 8134 8370 8186
rect 8422 8134 9292 8186
rect 1104 8112 9292 8134
rect 3234 8032 3240 8084
rect 3292 8032 3298 8084
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3375 8044 3801 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 5534 8032 5540 8084
rect 5592 8032 5598 8084
rect 5629 8075 5687 8081
rect 5629 8041 5641 8075
rect 5675 8072 5687 8075
rect 6914 8072 6920 8084
rect 5675 8044 6920 8072
rect 5675 8041 5687 8044
rect 5629 8035 5687 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 3050 8004 3056 8016
rect 2792 7976 3056 8004
rect 2792 7945 2820 7976
rect 3050 7964 3056 7976
rect 3108 8004 3114 8016
rect 3252 8004 3280 8032
rect 3421 8007 3479 8013
rect 3421 8004 3433 8007
rect 3108 7976 3280 8004
rect 3344 7976 3433 8004
rect 3108 7964 3114 7976
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3234 7868 3240 7880
rect 3007 7840 3240 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 2532 7803 2590 7809
rect 2532 7769 2544 7803
rect 2578 7800 2590 7803
rect 3344 7800 3372 7976
rect 3421 7973 3433 7976
rect 3467 7973 3479 8007
rect 3421 7967 3479 7973
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 7466 7936 7472 7948
rect 3568 7908 7472 7936
rect 3568 7896 3574 7908
rect 4080 7877 4108 7908
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 4065 7871 4123 7877
rect 3467 7840 3740 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 2578 7772 3372 7800
rect 2578 7769 2590 7772
rect 2532 7763 2590 7769
rect 1394 7692 1400 7744
rect 1452 7692 1458 7744
rect 2958 7692 2964 7744
rect 3016 7732 3022 7744
rect 3053 7735 3111 7741
rect 3053 7732 3065 7735
rect 3016 7704 3065 7732
rect 3016 7692 3022 7704
rect 3053 7701 3065 7704
rect 3099 7701 3111 7735
rect 3053 7695 3111 7701
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 3602 7732 3608 7744
rect 3191 7704 3608 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 3712 7732 3740 7840
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 9214 7868 9220 7880
rect 8711 7840 9220 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 3786 7760 3792 7812
rect 3844 7760 3850 7812
rect 3878 7760 3884 7812
rect 3936 7800 3942 7812
rect 3973 7803 4031 7809
rect 3973 7800 3985 7803
rect 3936 7772 3985 7800
rect 3936 7760 3942 7772
rect 3973 7769 3985 7772
rect 4019 7769 4031 7803
rect 5644 7800 5672 7831
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 5718 7800 5724 7812
rect 3973 7763 4031 7769
rect 5184 7772 5724 7800
rect 5184 7732 5212 7772
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 8478 7760 8484 7812
rect 8536 7760 8542 7812
rect 3712 7704 5212 7732
rect 5258 7692 5264 7744
rect 5316 7692 5322 7744
rect 5353 7735 5411 7741
rect 5353 7701 5365 7735
rect 5399 7732 5411 7735
rect 5442 7732 5448 7744
rect 5399 7704 5448 7732
rect 5399 7701 5411 7704
rect 5353 7695 5411 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 1104 7642 9292 7664
rect 1104 7590 2633 7642
rect 2685 7590 2697 7642
rect 2749 7590 2761 7642
rect 2813 7590 2825 7642
rect 2877 7590 2889 7642
rect 2941 7590 4680 7642
rect 4732 7590 4744 7642
rect 4796 7590 4808 7642
rect 4860 7590 4872 7642
rect 4924 7590 4936 7642
rect 4988 7590 6727 7642
rect 6779 7590 6791 7642
rect 6843 7590 6855 7642
rect 6907 7590 6919 7642
rect 6971 7590 6983 7642
rect 7035 7590 8774 7642
rect 8826 7590 8838 7642
rect 8890 7590 8902 7642
rect 8954 7590 8966 7642
rect 9018 7590 9030 7642
rect 9082 7590 9292 7642
rect 1104 7568 9292 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2958 7528 2964 7540
rect 2547 7500 2964 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3050 7488 3056 7540
rect 3108 7488 3114 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5316 7500 5365 7528
rect 5316 7488 5322 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5810 7528 5816 7540
rect 5353 7491 5411 7497
rect 5552 7500 5816 7528
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 2406 7460 2412 7472
rect 1636 7432 2176 7460
rect 1636 7420 1642 7432
rect 2148 7401 2176 7432
rect 2240 7432 2412 7460
rect 2240 7401 2268 7432
rect 2406 7420 2412 7432
rect 2464 7420 2470 7472
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 3326 7392 3332 7404
rect 2363 7364 3332 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2056 7324 2084 7355
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4338 7352 4344 7404
rect 4396 7352 4402 7404
rect 5552 7401 5580 7500
rect 5810 7488 5816 7500
rect 5868 7528 5874 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5868 7500 6377 7528
rect 5868 7488 5874 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6638 7420 6644 7472
rect 6696 7460 6702 7472
rect 7653 7463 7711 7469
rect 6696 7432 6776 7460
rect 6696 7420 6702 7432
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5629 7355 5687 7361
rect 5736 7364 5825 7392
rect 2056 7296 2360 7324
rect 2332 7200 2360 7296
rect 4430 7284 4436 7336
rect 4488 7324 4494 7336
rect 5258 7324 5264 7336
rect 4488 7296 5264 7324
rect 4488 7284 4494 7296
rect 5258 7284 5264 7296
rect 5316 7324 5322 7336
rect 5644 7324 5672 7355
rect 5316 7296 5672 7324
rect 5316 7284 5322 7296
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 5626 7256 5632 7268
rect 4672 7228 5632 7256
rect 4672 7216 4678 7228
rect 5626 7216 5632 7228
rect 5684 7256 5690 7268
rect 5736 7256 5764 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6748 7401 6776 7432
rect 7653 7429 7665 7463
rect 7699 7429 7711 7463
rect 7653 7423 7711 7429
rect 7869 7463 7927 7469
rect 7869 7429 7881 7463
rect 7915 7460 7927 7463
rect 8018 7460 8024 7472
rect 7915 7432 8024 7460
rect 7915 7429 7927 7432
rect 7869 7423 7927 7429
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 7668 7392 7696 7423
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 8662 7420 8668 7472
rect 8720 7420 8726 7472
rect 8680 7392 8708 7420
rect 7668 7364 8708 7392
rect 6733 7355 6791 7361
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 5684 7228 5764 7256
rect 5828 7296 6653 7324
rect 5684 7216 5690 7228
rect 5828 7200 5856 7296
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 2314 7148 2320 7200
rect 2372 7148 2378 7200
rect 5810 7148 5816 7200
rect 5868 7148 5874 7200
rect 7834 7148 7840 7200
rect 7892 7148 7898 7200
rect 7926 7148 7932 7200
rect 7984 7188 7990 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7984 7160 8033 7188
rect 7984 7148 7990 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 1104 7098 9292 7120
rect 1104 7046 1973 7098
rect 2025 7046 2037 7098
rect 2089 7046 2101 7098
rect 2153 7046 2165 7098
rect 2217 7046 2229 7098
rect 2281 7046 4020 7098
rect 4072 7046 4084 7098
rect 4136 7046 4148 7098
rect 4200 7046 4212 7098
rect 4264 7046 4276 7098
rect 4328 7046 6067 7098
rect 6119 7046 6131 7098
rect 6183 7046 6195 7098
rect 6247 7046 6259 7098
rect 6311 7046 6323 7098
rect 6375 7046 8114 7098
rect 8166 7046 8178 7098
rect 8230 7046 8242 7098
rect 8294 7046 8306 7098
rect 8358 7046 8370 7098
rect 8422 7046 9292 7098
rect 1104 7024 9292 7046
rect 3234 6944 3240 6996
rect 3292 6944 3298 6996
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 5442 6984 5448 6996
rect 3844 6956 5448 6984
rect 3844 6944 3850 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 5534 6944 5540 6996
rect 5592 6944 5598 6996
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 5994 6984 6000 6996
rect 5776 6956 6000 6984
rect 5776 6944 5782 6956
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7892 6956 8125 6984
rect 7892 6944 7898 6956
rect 8113 6953 8125 6956
rect 8159 6953 8171 6987
rect 8113 6947 8171 6953
rect 5902 6916 5908 6928
rect 1596 6888 5908 6916
rect 1596 6860 1624 6888
rect 1578 6808 1584 6860
rect 1636 6808 1642 6860
rect 3142 6848 3148 6860
rect 2976 6820 3148 6848
rect 2976 6789 3004 6820
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 4473 6857 4501 6888
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 7926 6916 7932 6928
rect 7392 6888 7932 6916
rect 4458 6851 4516 6857
rect 4458 6817 4470 6851
rect 4504 6817 4516 6851
rect 4458 6811 4516 6817
rect 4614 6808 4620 6860
rect 4672 6808 4678 6860
rect 7392 6857 7420 6888
rect 7926 6876 7932 6888
rect 7984 6876 7990 6928
rect 7377 6851 7435 6857
rect 5736 6820 6684 6848
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3108 6752 3985 6780
rect 3108 6740 3114 6752
rect 3973 6749 3985 6752
rect 4019 6780 4031 6783
rect 4632 6780 4660 6808
rect 5736 6792 5764 6820
rect 6656 6792 6684 6820
rect 7377 6817 7389 6851
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 7466 6808 7472 6860
rect 7524 6808 7530 6860
rect 7760 6820 7972 6848
rect 4019 6752 4660 6780
rect 4019 6749 4031 6752
rect 3973 6743 4031 6749
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 3234 6672 3240 6724
rect 3292 6672 3298 6724
rect 3418 6672 3424 6724
rect 3476 6712 3482 6724
rect 4341 6715 4399 6721
rect 4341 6712 4353 6715
rect 3476 6684 4353 6712
rect 3476 6672 3482 6684
rect 4341 6681 4353 6684
rect 4387 6712 4399 6715
rect 4430 6712 4436 6724
rect 4387 6684 4436 6712
rect 4387 6681 4399 6684
rect 4341 6675 4399 6681
rect 4430 6672 4436 6684
rect 4488 6672 4494 6724
rect 5534 6672 5540 6724
rect 5592 6672 5598 6724
rect 5828 6656 5856 6743
rect 6638 6740 6644 6792
rect 6696 6740 6702 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 7147 6783 7205 6789
rect 7147 6749 7159 6783
rect 7193 6780 7205 6783
rect 7650 6780 7656 6792
rect 7193 6752 7656 6780
rect 7193 6749 7205 6752
rect 7147 6743 7205 6749
rect 7024 6712 7052 6743
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 7760 6724 7788 6820
rect 7944 6789 7972 6820
rect 8018 6808 8024 6860
rect 8076 6808 8082 6860
rect 8128 6848 8156 6947
rect 8128 6820 8340 6848
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 8036 6780 8064 6808
rect 8312 6789 8340 6820
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 8036 6752 8217 6780
rect 7929 6743 7987 6749
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6780 8539 6783
rect 8662 6780 8668 6792
rect 8527 6752 8668 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 7558 6712 7564 6724
rect 7024 6684 7564 6712
rect 7558 6672 7564 6684
rect 7616 6672 7622 6724
rect 7742 6672 7748 6724
rect 7800 6672 7806 6724
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3602 6644 3608 6656
rect 3099 6616 3608 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 4246 6644 4252 6656
rect 3844 6616 4252 6644
rect 3844 6604 3850 6616
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 5074 6644 5080 6656
rect 4663 6616 5080 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5810 6604 5816 6656
rect 5868 6604 5874 6656
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6644 7067 6647
rect 7098 6644 7104 6656
rect 7055 6616 7104 6644
rect 7055 6613 7067 6616
rect 7009 6607 7067 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7852 6644 7880 6743
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 7340 6616 7880 6644
rect 7340 6604 7346 6616
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 8628 6616 8677 6644
rect 8628 6604 8634 6616
rect 8665 6613 8677 6616
rect 8711 6613 8723 6647
rect 8665 6607 8723 6613
rect 1104 6554 9292 6576
rect 1104 6502 2633 6554
rect 2685 6502 2697 6554
rect 2749 6502 2761 6554
rect 2813 6502 2825 6554
rect 2877 6502 2889 6554
rect 2941 6502 4680 6554
rect 4732 6502 4744 6554
rect 4796 6502 4808 6554
rect 4860 6502 4872 6554
rect 4924 6502 4936 6554
rect 4988 6502 6727 6554
rect 6779 6502 6791 6554
rect 6843 6502 6855 6554
rect 6907 6502 6919 6554
rect 6971 6502 6983 6554
rect 7035 6502 8774 6554
rect 8826 6502 8838 6554
rect 8890 6502 8902 6554
rect 8954 6502 8966 6554
rect 9018 6502 9030 6554
rect 9082 6502 9292 6554
rect 1104 6480 9292 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 2314 6440 2320 6452
rect 1811 6412 2320 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 2314 6400 2320 6412
rect 2372 6440 2378 6452
rect 2803 6443 2861 6449
rect 2803 6440 2815 6443
rect 2372 6412 2815 6440
rect 2372 6400 2378 6412
rect 2803 6409 2815 6412
rect 2849 6440 2861 6443
rect 3050 6440 3056 6452
rect 2849 6412 3056 6440
rect 2849 6409 2861 6412
rect 2803 6403 2861 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 3292 6412 3709 6440
rect 3292 6400 3298 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 4801 6443 4859 6449
rect 4801 6440 4813 6443
rect 3697 6403 3755 6409
rect 3988 6412 4813 6440
rect 2041 6375 2099 6381
rect 2041 6341 2053 6375
rect 2087 6372 2099 6375
rect 2406 6372 2412 6384
rect 2087 6344 2412 6372
rect 2087 6341 2099 6344
rect 2041 6335 2099 6341
rect 2406 6332 2412 6344
rect 2464 6372 2470 6384
rect 2593 6375 2651 6381
rect 2593 6372 2605 6375
rect 2464 6344 2605 6372
rect 2464 6332 2470 6344
rect 2593 6341 2605 6344
rect 2639 6372 2651 6375
rect 3418 6372 3424 6384
rect 2639 6344 3424 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 3418 6332 3424 6344
rect 3476 6332 3482 6384
rect 3988 6381 4016 6412
rect 4801 6409 4813 6412
rect 4847 6440 4859 6443
rect 4847 6412 5764 6440
rect 4847 6409 4859 6412
rect 4801 6403 4859 6409
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6341 4031 6375
rect 3973 6335 4031 6341
rect 5074 6332 5080 6384
rect 5132 6332 5138 6384
rect 5166 6332 5172 6384
rect 5224 6332 5230 6384
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 3878 6313 3884 6316
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1912 6276 1961 6304
rect 1912 6264 1918 6276
rect 1949 6273 1961 6276
rect 1995 6304 2007 6307
rect 3876 6304 3884 6313
rect 1995 6276 2452 6304
rect 3839 6276 3884 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2314 6128 2320 6180
rect 2372 6128 2378 6180
rect 2424 6168 2452 6276
rect 3876 6267 3884 6276
rect 3878 6264 3884 6267
rect 3936 6264 3942 6316
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6273 4123 6307
rect 4246 6304 4252 6316
rect 4207 6276 4252 6304
rect 4065 6267 4123 6273
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 3602 6236 3608 6248
rect 2547 6208 3608 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 4080 6236 4108 6267
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 4522 6304 4528 6316
rect 4387 6276 4528 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5092 6304 5120 6332
rect 5736 6316 5764 6412
rect 7558 6400 7564 6452
rect 7616 6440 7622 6452
rect 7616 6412 7972 6440
rect 7616 6400 7622 6412
rect 7282 6332 7288 6384
rect 7340 6372 7346 6384
rect 7340 6344 7788 6372
rect 7340 6332 7346 6344
rect 5031 6276 5120 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 4724 6236 4752 6267
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 7760 6313 7788 6344
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7524 6276 7665 6304
rect 7524 6264 7530 6276
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 7834 6264 7840 6316
rect 7892 6264 7898 6316
rect 7944 6304 7972 6412
rect 8018 6400 8024 6452
rect 8076 6400 8082 6452
rect 8570 6304 8576 6316
rect 7944 6276 8576 6304
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 4080 6208 4752 6236
rect 2961 6171 3019 6177
rect 2424 6140 2912 6168
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 1854 6100 1860 6112
rect 1636 6072 1860 6100
rect 1636 6060 1642 6072
rect 1854 6060 1860 6072
rect 1912 6100 1918 6112
rect 2777 6103 2835 6109
rect 2777 6100 2789 6103
rect 1912 6072 2789 6100
rect 1912 6060 1918 6072
rect 2777 6069 2789 6072
rect 2823 6069 2835 6103
rect 2884 6100 2912 6140
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 3050 6168 3056 6180
rect 3007 6140 3056 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 3050 6128 3056 6140
rect 3108 6168 3114 6180
rect 4080 6168 4108 6208
rect 3108 6140 4108 6168
rect 4724 6168 4752 6208
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5123 6208 5273 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5261 6205 5273 6208
rect 5307 6205 5319 6239
rect 5261 6199 5319 6205
rect 5166 6168 5172 6180
rect 4724 6140 5172 6168
rect 3108 6128 3114 6140
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 5718 6128 5724 6180
rect 5776 6168 5782 6180
rect 5994 6168 6000 6180
rect 5776 6140 6000 6168
rect 5776 6128 5782 6140
rect 5994 6128 6000 6140
rect 6052 6128 6058 6180
rect 7926 6128 7932 6180
rect 7984 6168 7990 6180
rect 8113 6171 8171 6177
rect 8113 6168 8125 6171
rect 7984 6140 8125 6168
rect 7984 6128 7990 6140
rect 8113 6137 8125 6140
rect 8159 6137 8171 6171
rect 8113 6131 8171 6137
rect 5534 6100 5540 6112
rect 2884 6072 5540 6100
rect 2777 6063 2835 6069
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 5810 6100 5816 6112
rect 5675 6072 5816 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 5810 6060 5816 6072
rect 5868 6100 5874 6112
rect 7742 6100 7748 6112
rect 5868 6072 7748 6100
rect 5868 6060 5874 6072
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 8297 6103 8355 6109
rect 8297 6100 8309 6103
rect 8076 6072 8309 6100
rect 8076 6060 8082 6072
rect 8297 6069 8309 6072
rect 8343 6069 8355 6103
rect 8297 6063 8355 6069
rect 1104 6010 9292 6032
rect 1104 5958 1973 6010
rect 2025 5958 2037 6010
rect 2089 5958 2101 6010
rect 2153 5958 2165 6010
rect 2217 5958 2229 6010
rect 2281 5958 4020 6010
rect 4072 5958 4084 6010
rect 4136 5958 4148 6010
rect 4200 5958 4212 6010
rect 4264 5958 4276 6010
rect 4328 5958 6067 6010
rect 6119 5958 6131 6010
rect 6183 5958 6195 6010
rect 6247 5958 6259 6010
rect 6311 5958 6323 6010
rect 6375 5958 8114 6010
rect 8166 5958 8178 6010
rect 8230 5958 8242 6010
rect 8294 5958 8306 6010
rect 8358 5958 8370 6010
rect 8422 5958 9292 6010
rect 1104 5936 9292 5958
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4522 5896 4528 5908
rect 4387 5868 4528 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 5920 5868 7420 5896
rect 5920 5840 5948 5868
rect 4433 5831 4491 5837
rect 4433 5797 4445 5831
rect 4479 5797 4491 5831
rect 4433 5791 4491 5797
rect 4985 5831 5043 5837
rect 4985 5797 4997 5831
rect 5031 5828 5043 5831
rect 5258 5828 5264 5840
rect 5031 5800 5264 5828
rect 5031 5797 5043 5800
rect 4985 5791 5043 5797
rect 3510 5720 3516 5772
rect 3568 5760 3574 5772
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 3568 5732 3893 5760
rect 3568 5720 3574 5732
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 4448 5760 4476 5791
rect 5258 5788 5264 5800
rect 5316 5788 5322 5840
rect 5902 5788 5908 5840
rect 5960 5788 5966 5840
rect 6546 5788 6552 5840
rect 6604 5788 6610 5840
rect 3881 5723 3939 5729
rect 4080 5732 4476 5760
rect 5552 5732 7328 5760
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1489 5695 1547 5701
rect 1489 5692 1501 5695
rect 1452 5664 1501 5692
rect 1452 5652 1458 5664
rect 1489 5661 1501 5664
rect 1535 5661 1547 5695
rect 1489 5655 1547 5661
rect 2958 5652 2964 5704
rect 3016 5692 3022 5704
rect 3786 5692 3792 5704
rect 3016 5664 3792 5692
rect 3016 5652 3022 5664
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 3804 5556 3832 5652
rect 3896 5624 3924 5723
rect 4080 5701 4108 5732
rect 5552 5704 5580 5732
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 4423 5695 4481 5701
rect 4423 5661 4435 5695
rect 4469 5692 4481 5695
rect 4614 5692 4620 5704
rect 4469 5664 4620 5692
rect 4469 5661 4481 5664
rect 4423 5655 4481 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 4724 5624 4752 5655
rect 3896 5596 4752 5624
rect 4617 5559 4675 5565
rect 4617 5556 4629 5559
rect 3804 5528 4629 5556
rect 4617 5525 4629 5528
rect 4663 5525 4675 5559
rect 5184 5556 5212 5655
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 7300 5701 7328 5732
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5661 7343 5695
rect 7392 5692 7420 5868
rect 7834 5788 7840 5840
rect 7892 5788 7898 5840
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7392 5664 7481 5692
rect 7285 5655 7343 5661
rect 7469 5661 7481 5664
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 8803 5664 9352 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 5258 5584 5264 5636
rect 5316 5584 5322 5636
rect 6638 5556 6644 5568
rect 5184 5528 6644 5556
rect 4617 5519 4675 5525
rect 6638 5516 6644 5528
rect 6696 5556 6702 5568
rect 7208 5556 7236 5655
rect 9324 5568 9352 5664
rect 8573 5559 8631 5565
rect 8573 5556 8585 5559
rect 6696 5528 8585 5556
rect 6696 5516 6702 5528
rect 8573 5525 8585 5528
rect 8619 5525 8631 5559
rect 8573 5519 8631 5525
rect 9306 5516 9312 5568
rect 9364 5516 9370 5568
rect 1104 5466 9292 5488
rect 1104 5414 2633 5466
rect 2685 5414 2697 5466
rect 2749 5414 2761 5466
rect 2813 5414 2825 5466
rect 2877 5414 2889 5466
rect 2941 5414 4680 5466
rect 4732 5414 4744 5466
rect 4796 5414 4808 5466
rect 4860 5414 4872 5466
rect 4924 5414 4936 5466
rect 4988 5414 6727 5466
rect 6779 5414 6791 5466
rect 6843 5414 6855 5466
rect 6907 5414 6919 5466
rect 6971 5414 6983 5466
rect 7035 5414 8774 5466
rect 8826 5414 8838 5466
rect 8890 5414 8902 5466
rect 8954 5414 8966 5466
rect 9018 5414 9030 5466
rect 9082 5414 9292 5466
rect 1104 5392 9292 5414
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5352 2283 5355
rect 2406 5352 2412 5364
rect 2271 5324 2412 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 2685 5355 2743 5361
rect 2685 5321 2697 5355
rect 2731 5321 2743 5355
rect 2685 5315 2743 5321
rect 2700 5284 2728 5315
rect 3602 5312 3608 5364
rect 3660 5312 3666 5364
rect 3786 5312 3792 5364
rect 3844 5352 3850 5364
rect 4154 5352 4160 5364
rect 3844 5324 4160 5352
rect 3844 5312 3850 5324
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 4488 5324 5641 5352
rect 4488 5312 4494 5324
rect 5629 5321 5641 5324
rect 5675 5321 5687 5355
rect 5629 5315 5687 5321
rect 7558 5312 7564 5364
rect 7616 5312 7622 5364
rect 3421 5287 3479 5293
rect 3421 5284 3433 5287
rect 2700 5256 3433 5284
rect 3421 5253 3433 5256
rect 3467 5253 3479 5287
rect 5074 5284 5080 5296
rect 3421 5247 3479 5253
rect 5000 5256 5080 5284
rect 1854 5176 1860 5228
rect 1912 5176 1918 5228
rect 2864 5219 2922 5225
rect 2864 5185 2876 5219
rect 2910 5185 2922 5219
rect 2864 5179 2922 5185
rect 2879 5148 2907 5179
rect 2958 5176 2964 5228
rect 3016 5176 3022 5228
rect 3050 5176 3056 5228
rect 3108 5176 3114 5228
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3326 5176 3332 5228
rect 3384 5176 3390 5228
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 4890 5216 4896 5228
rect 3743 5188 4896 5216
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 5000 5225 5028 5256
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 5166 5244 5172 5296
rect 5224 5244 5230 5296
rect 5261 5287 5319 5293
rect 5261 5253 5273 5287
rect 5307 5284 5319 5287
rect 5307 5256 5488 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 5460 5228 5488 5256
rect 7852 5256 8708 5284
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 5353 5219 5411 5225
rect 5353 5206 5365 5219
rect 4985 5179 5043 5185
rect 5092 5185 5365 5206
rect 5399 5185 5411 5219
rect 5092 5179 5411 5185
rect 5092 5178 5396 5179
rect 3878 5148 3884 5160
rect 2879 5120 3884 5148
rect 2409 5083 2467 5089
rect 2409 5049 2421 5083
rect 2455 5080 2467 5083
rect 2879 5080 2907 5120
rect 3878 5108 3884 5120
rect 3936 5148 3942 5160
rect 5092 5148 5120 5178
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 5534 5176 5540 5228
rect 5592 5176 5598 5228
rect 5902 5176 5908 5228
rect 5960 5176 5966 5228
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6638 5216 6644 5228
rect 6227 5188 6644 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 7852 5216 7880 5256
rect 7340 5188 7880 5216
rect 7340 5176 7346 5188
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8680 5225 8708 5256
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 3936 5120 5120 5148
rect 3936 5108 3942 5120
rect 2455 5052 2907 5080
rect 5552 5080 5580 5176
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 7708 5120 7849 5148
rect 7708 5108 7714 5120
rect 7837 5117 7849 5120
rect 7883 5148 7895 5151
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7883 5120 8217 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 5552 5052 5856 5080
rect 2455 5049 2467 5052
rect 2409 5043 2467 5049
rect 2225 5015 2283 5021
rect 2225 4981 2237 5015
rect 2271 5012 2283 5015
rect 2314 5012 2320 5024
rect 2271 4984 2320 5012
rect 2271 4981 2283 4984
rect 2225 4975 2283 4981
rect 2314 4972 2320 4984
rect 2372 4972 2378 5024
rect 3418 4972 3424 5024
rect 3476 4972 3482 5024
rect 5534 4972 5540 5024
rect 5592 4972 5598 5024
rect 5828 5021 5856 5052
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 4981 5871 5015
rect 5813 4975 5871 4981
rect 8478 4972 8484 5024
rect 8536 4972 8542 5024
rect 1104 4922 9292 4944
rect 1104 4870 1973 4922
rect 2025 4870 2037 4922
rect 2089 4870 2101 4922
rect 2153 4870 2165 4922
rect 2217 4870 2229 4922
rect 2281 4870 4020 4922
rect 4072 4870 4084 4922
rect 4136 4870 4148 4922
rect 4200 4870 4212 4922
rect 4264 4870 4276 4922
rect 4328 4870 6067 4922
rect 6119 4870 6131 4922
rect 6183 4870 6195 4922
rect 6247 4870 6259 4922
rect 6311 4870 6323 4922
rect 6375 4870 8114 4922
rect 8166 4870 8178 4922
rect 8230 4870 8242 4922
rect 8294 4870 8306 4922
rect 8358 4870 8370 4922
rect 8422 4870 9292 4922
rect 1104 4848 9292 4870
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3384 4780 3801 4808
rect 3384 4768 3390 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5408 4780 5825 4808
rect 5408 4768 5414 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 6454 4808 6460 4820
rect 6227 4780 6460 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 4433 4743 4491 4749
rect 4433 4740 4445 4743
rect 4080 4712 4445 4740
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4080 4613 4108 4712
rect 4433 4709 4445 4712
rect 4479 4709 4491 4743
rect 4433 4703 4491 4709
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4522 4672 4528 4684
rect 4295 4644 4528 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4522 4632 4528 4644
rect 4580 4672 4586 4684
rect 4580 4644 4752 4672
rect 4580 4632 4586 4644
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 3234 4496 3240 4548
rect 3292 4536 3298 4548
rect 4356 4536 4384 4567
rect 4430 4564 4436 4616
rect 4488 4564 4494 4616
rect 4724 4613 4752 4644
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 5644 4604 5672 4700
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5644 4576 5733 4604
rect 4709 4567 4767 4573
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 4724 4536 4752 4567
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 7484 4536 7512 4564
rect 3292 4508 4660 4536
rect 4724 4508 7512 4536
rect 3292 4496 3298 4508
rect 4632 4477 4660 4508
rect 8662 4496 8668 4548
rect 8720 4496 8726 4548
rect 4617 4471 4675 4477
rect 4617 4437 4629 4471
rect 4663 4468 4675 4471
rect 5166 4468 5172 4480
rect 4663 4440 5172 4468
rect 4663 4437 4675 4440
rect 4617 4431 4675 4437
rect 5166 4428 5172 4440
rect 5224 4468 5230 4480
rect 5442 4468 5448 4480
rect 5224 4440 5448 4468
rect 5224 4428 5230 4440
rect 5442 4428 5448 4440
rect 5500 4468 5506 4480
rect 8680 4468 8708 4496
rect 5500 4440 8708 4468
rect 5500 4428 5506 4440
rect 1104 4378 9292 4400
rect 1104 4326 2633 4378
rect 2685 4326 2697 4378
rect 2749 4326 2761 4378
rect 2813 4326 2825 4378
rect 2877 4326 2889 4378
rect 2941 4326 4680 4378
rect 4732 4326 4744 4378
rect 4796 4326 4808 4378
rect 4860 4326 4872 4378
rect 4924 4326 4936 4378
rect 4988 4326 6727 4378
rect 6779 4326 6791 4378
rect 6843 4326 6855 4378
rect 6907 4326 6919 4378
rect 6971 4326 6983 4378
rect 7035 4326 8774 4378
rect 8826 4326 8838 4378
rect 8890 4326 8902 4378
rect 8954 4326 8966 4378
rect 9018 4326 9030 4378
rect 9082 4326 9292 4378
rect 1104 4304 9292 4326
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 6638 4264 6644 4276
rect 5868 4236 6644 4264
rect 5868 4224 5874 4236
rect 6638 4224 6644 4236
rect 6696 4264 6702 4276
rect 6696 4236 6960 4264
rect 6696 4224 6702 4236
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 5721 4199 5779 4205
rect 5721 4196 5733 4199
rect 4488 4168 5733 4196
rect 4488 4156 4494 4168
rect 5721 4165 5733 4168
rect 5767 4165 5779 4199
rect 5721 4159 5779 4165
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 5828 4128 5856 4224
rect 5905 4199 5963 4205
rect 5905 4165 5917 4199
rect 5951 4196 5963 4199
rect 6454 4196 6460 4208
rect 5951 4168 6460 4196
rect 5951 4165 5963 4168
rect 5905 4159 5963 4165
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6564 4168 6776 4196
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 3936 4100 6009 4128
rect 3936 4088 3942 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6125 4131 6183 4137
rect 6125 4097 6137 4131
rect 6171 4128 6183 4131
rect 6362 4128 6368 4140
rect 6171 4100 6368 4128
rect 6171 4097 6183 4100
rect 6125 4091 6183 4097
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6564 4137 6592 4168
rect 6550 4131 6608 4137
rect 6550 4097 6562 4131
rect 6596 4097 6608 4131
rect 6550 4091 6608 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 5905 4063 5963 4069
rect 5905 4029 5917 4063
rect 5951 4060 5963 4063
rect 6656 4060 6684 4091
rect 5951 4032 6684 4060
rect 5951 4029 5963 4032
rect 5905 4023 5963 4029
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 5166 3992 5172 4004
rect 4028 3964 5172 3992
rect 4028 3952 4034 3964
rect 5166 3952 5172 3964
rect 5224 3992 5230 4004
rect 6748 3992 6776 4168
rect 6932 4137 6960 4236
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 8478 4128 8484 4140
rect 6963 4100 8484 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7282 4060 7288 4072
rect 6871 4032 7288 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 5224 3964 6776 3992
rect 5224 3952 5230 3964
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5960 3896 6377 3924
rect 5960 3884 5966 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 6840 3924 6868 4023
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 6512 3896 6868 3924
rect 6512 3884 6518 3896
rect 1104 3834 9292 3856
rect 1104 3782 1973 3834
rect 2025 3782 2037 3834
rect 2089 3782 2101 3834
rect 2153 3782 2165 3834
rect 2217 3782 2229 3834
rect 2281 3782 4020 3834
rect 4072 3782 4084 3834
rect 4136 3782 4148 3834
rect 4200 3782 4212 3834
rect 4264 3782 4276 3834
rect 4328 3782 6067 3834
rect 6119 3782 6131 3834
rect 6183 3782 6195 3834
rect 6247 3782 6259 3834
rect 6311 3782 6323 3834
rect 6375 3782 8114 3834
rect 8166 3782 8178 3834
rect 8230 3782 8242 3834
rect 8294 3782 8306 3834
rect 8358 3782 8370 3834
rect 8422 3782 9292 3834
rect 1104 3760 9292 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 2409 3723 2467 3729
rect 2409 3720 2421 3723
rect 1912 3692 2421 3720
rect 1912 3680 1918 3692
rect 2409 3689 2421 3692
rect 2455 3689 2467 3723
rect 2409 3683 2467 3689
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 3694 3720 3700 3732
rect 3283 3692 3700 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 2314 3612 2320 3664
rect 2372 3612 2378 3664
rect 2332 3516 2360 3612
rect 2424 3584 2452 3683
rect 3694 3680 3700 3692
rect 3752 3720 3758 3732
rect 3752 3692 5488 3720
rect 3752 3680 3758 3692
rect 2608 3624 5304 3652
rect 2424 3556 2544 3584
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 2332 3488 2421 3516
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 1486 3408 1492 3460
rect 1544 3408 1550 3460
rect 2516 3448 2544 3556
rect 2608 3525 2636 3624
rect 4080 3525 4108 3624
rect 4356 3556 4844 3584
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 2593 3479 2651 3485
rect 2700 3488 3985 3516
rect 2700 3448 2728 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 3145 3451 3203 3457
rect 3145 3448 3157 3451
rect 2516 3420 2728 3448
rect 2792 3420 3157 3448
rect 934 3340 940 3392
rect 992 3380 998 3392
rect 2792 3389 2820 3420
rect 3145 3417 3157 3420
rect 3191 3417 3203 3451
rect 3988 3448 4016 3479
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4267 3519 4325 3525
rect 4267 3485 4279 3519
rect 4313 3516 4325 3519
rect 4356 3516 4384 3556
rect 4816 3525 4844 3556
rect 5276 3525 5304 3624
rect 4313 3488 4384 3516
rect 4433 3519 4491 3525
rect 4313 3485 4325 3488
rect 4267 3479 4325 3485
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5350 3516 5356 3528
rect 5307 3488 5356 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 4448 3448 4476 3479
rect 3988 3420 4476 3448
rect 4816 3448 4844 3479
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5460 3516 5488 3692
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5592 3692 5641 3720
rect 5592 3680 5598 3692
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 5629 3683 5687 3689
rect 5902 3680 5908 3732
rect 5960 3680 5966 3732
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 5920 3584 5948 3680
rect 5859 3556 5948 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 5460 3488 5549 3516
rect 5537 3485 5549 3488
rect 5583 3516 5595 3519
rect 6546 3516 6552 3528
rect 5583 3488 6552 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 5626 3448 5632 3460
rect 4816 3420 5632 3448
rect 3145 3411 3203 3417
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 992 3352 1593 3380
rect 992 3340 998 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 2777 3383 2835 3389
rect 2777 3349 2789 3383
rect 2823 3349 2835 3383
rect 2777 3343 2835 3349
rect 3786 3340 3792 3392
rect 3844 3340 3850 3392
rect 5166 3340 5172 3392
rect 5224 3340 5230 3392
rect 5902 3340 5908 3392
rect 5960 3380 5966 3392
rect 6089 3383 6147 3389
rect 6089 3380 6101 3383
rect 5960 3352 6101 3380
rect 5960 3340 5966 3352
rect 6089 3349 6101 3352
rect 6135 3349 6147 3383
rect 6089 3343 6147 3349
rect 1104 3290 9292 3312
rect 1104 3238 2633 3290
rect 2685 3238 2697 3290
rect 2749 3238 2761 3290
rect 2813 3238 2825 3290
rect 2877 3238 2889 3290
rect 2941 3238 4680 3290
rect 4732 3238 4744 3290
rect 4796 3238 4808 3290
rect 4860 3238 4872 3290
rect 4924 3238 4936 3290
rect 4988 3238 6727 3290
rect 6779 3238 6791 3290
rect 6843 3238 6855 3290
rect 6907 3238 6919 3290
rect 6971 3238 6983 3290
rect 7035 3238 8774 3290
rect 8826 3238 8838 3290
rect 8890 3238 8902 3290
rect 8954 3238 8966 3290
rect 9018 3238 9030 3290
rect 9082 3238 9292 3290
rect 1104 3216 9292 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 4522 3176 4528 3188
rect 1627 3148 4528 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 5074 3176 5080 3188
rect 4663 3148 5080 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 6454 3136 6460 3188
rect 6512 3136 6518 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 6733 3179 6791 3185
rect 6733 3176 6745 3179
rect 6696 3148 6745 3176
rect 6696 3136 6702 3148
rect 6733 3145 6745 3148
rect 6779 3145 6791 3179
rect 6733 3139 6791 3145
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 8573 3179 8631 3185
rect 8573 3145 8585 3179
rect 8619 3145 8631 3179
rect 8573 3139 8631 3145
rect 3694 3068 3700 3120
rect 3752 3068 3758 3120
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 14 3000 20 3052
rect 72 3040 78 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 72 3012 1501 3040
rect 72 3000 78 3012
rect 1489 3009 1501 3012
rect 1535 3009 1547 3043
rect 3712 3040 3740 3068
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 3712 3012 4445 3040
rect 1489 3003 1547 3009
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4540 3040 4568 3136
rect 5905 3111 5963 3117
rect 5905 3077 5917 3111
rect 5951 3108 5963 3111
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 5951 3080 6377 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 6472 3108 6500 3136
rect 7116 3108 7144 3139
rect 7438 3111 7496 3117
rect 7438 3108 7450 3111
rect 6472 3080 6684 3108
rect 7116 3080 7450 3108
rect 6365 3071 6423 3077
rect 4709 3043 4767 3049
rect 4709 3040 4721 3043
rect 4540 3012 4721 3040
rect 4433 3003 4491 3009
rect 4709 3009 4721 3012
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5718 3040 5724 3052
rect 5583 3012 5724 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 6656 3040 6684 3080
rect 7438 3077 7450 3080
rect 7484 3077 7496 3111
rect 7438 3071 7496 3077
rect 6825 3044 6883 3049
rect 6748 3043 6883 3044
rect 6748 3040 6837 3043
rect 6656 3016 6837 3040
rect 6656 3012 6776 3016
rect 6825 3009 6837 3016
rect 6871 3009 6883 3043
rect 7193 3043 7251 3049
rect 6825 3003 6883 3009
rect 6917 3027 6975 3033
rect 6917 2993 6929 3027
rect 6963 3024 6975 3027
rect 6963 2996 7052 3024
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 8588 3040 8616 3139
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8588 3012 8677 3040
rect 7193 3003 7251 3009
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 6963 2993 6975 2996
rect 6917 2987 6975 2993
rect 3068 2944 6040 2972
rect 3068 2916 3096 2944
rect 3050 2864 3056 2916
rect 3108 2864 3114 2916
rect 4430 2796 4436 2848
rect 4488 2796 4494 2848
rect 5902 2796 5908 2848
rect 5960 2796 5966 2848
rect 6012 2836 6040 2944
rect 6089 2907 6147 2913
rect 6089 2873 6101 2907
rect 6135 2904 6147 2907
rect 7024 2904 7052 2996
rect 6135 2876 7052 2904
rect 6135 2873 6147 2876
rect 6089 2867 6147 2873
rect 7208 2836 7236 3003
rect 6012 2808 7236 2836
rect 8846 2796 8852 2848
rect 8904 2796 8910 2848
rect 1104 2746 9292 2768
rect 1104 2694 1973 2746
rect 2025 2694 2037 2746
rect 2089 2694 2101 2746
rect 2153 2694 2165 2746
rect 2217 2694 2229 2746
rect 2281 2694 4020 2746
rect 4072 2694 4084 2746
rect 4136 2694 4148 2746
rect 4200 2694 4212 2746
rect 4264 2694 4276 2746
rect 4328 2694 6067 2746
rect 6119 2694 6131 2746
rect 6183 2694 6195 2746
rect 6247 2694 6259 2746
rect 6311 2694 6323 2746
rect 6375 2694 8114 2746
rect 8166 2694 8178 2746
rect 8230 2694 8242 2746
rect 8294 2694 8306 2746
rect 8358 2694 8370 2746
rect 8422 2694 9292 2746
rect 1104 2672 9292 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 1486 2632 1492 2644
rect 1443 2604 1492 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 1486 2592 1492 2604
rect 1544 2592 1550 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4430 2632 4436 2644
rect 4203 2604 4436 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5626 2632 5632 2644
rect 5491 2604 5632 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3050 2496 3056 2508
rect 2823 2468 3056 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 5460 2496 5488 2595
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 7834 2592 7840 2644
rect 7892 2592 7898 2644
rect 8573 2635 8631 2641
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 8662 2632 8668 2644
rect 8619 2604 8668 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 4264 2468 5488 2496
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3476 2400 3801 2428
rect 3476 2388 3482 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3878 2388 3884 2440
rect 3936 2388 3942 2440
rect 4264 2437 4292 2468
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 10318 2428 10324 2440
rect 8803 2400 10324 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 2532 2363 2590 2369
rect 2532 2329 2544 2363
rect 2578 2360 2590 2363
rect 2578 2332 4292 2360
rect 2578 2329 2590 2332
rect 2532 2323 2590 2329
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 4264 2301 4292 2332
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3568 2264 3985 2292
rect 3568 2252 3574 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 4249 2295 4307 2301
rect 4249 2261 4261 2295
rect 4295 2261 4307 2295
rect 4249 2255 4307 2261
rect 1104 2202 9292 2224
rect 1104 2150 2633 2202
rect 2685 2150 2697 2202
rect 2749 2150 2761 2202
rect 2813 2150 2825 2202
rect 2877 2150 2889 2202
rect 2941 2150 4680 2202
rect 4732 2150 4744 2202
rect 4796 2150 4808 2202
rect 4860 2150 4872 2202
rect 4924 2150 4936 2202
rect 4988 2150 6727 2202
rect 6779 2150 6791 2202
rect 6843 2150 6855 2202
rect 6907 2150 6919 2202
rect 6971 2150 6983 2202
rect 7035 2150 8774 2202
rect 8826 2150 8838 2202
rect 8890 2150 8902 2202
rect 8954 2150 8966 2202
rect 9018 2150 9030 2202
rect 9082 2150 9292 2202
rect 1104 2128 9292 2150
<< via1 >>
rect 1973 10310 2025 10362
rect 2037 10310 2089 10362
rect 2101 10310 2153 10362
rect 2165 10310 2217 10362
rect 2229 10310 2281 10362
rect 4020 10310 4072 10362
rect 4084 10310 4136 10362
rect 4148 10310 4200 10362
rect 4212 10310 4264 10362
rect 4276 10310 4328 10362
rect 6067 10310 6119 10362
rect 6131 10310 6183 10362
rect 6195 10310 6247 10362
rect 6259 10310 6311 10362
rect 6323 10310 6375 10362
rect 8114 10310 8166 10362
rect 8178 10310 8230 10362
rect 8242 10310 8294 10362
rect 8306 10310 8358 10362
rect 8370 10310 8422 10362
rect 1308 10208 1360 10260
rect 9036 10208 9088 10260
rect 2964 10140 3016 10192
rect 940 10004 992 10056
rect 3884 10004 3936 10056
rect 6460 10004 6512 10056
rect 9220 10004 9272 10056
rect 7104 9936 7156 9988
rect 8484 9936 8536 9988
rect 1860 9868 1912 9920
rect 6644 9868 6696 9920
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 2633 9766 2685 9818
rect 2697 9766 2749 9818
rect 2761 9766 2813 9818
rect 2825 9766 2877 9818
rect 2889 9766 2941 9818
rect 4680 9766 4732 9818
rect 4744 9766 4796 9818
rect 4808 9766 4860 9818
rect 4872 9766 4924 9818
rect 4936 9766 4988 9818
rect 6727 9766 6779 9818
rect 6791 9766 6843 9818
rect 6855 9766 6907 9818
rect 6919 9766 6971 9818
rect 6983 9766 7035 9818
rect 8774 9766 8826 9818
rect 8838 9766 8890 9818
rect 8902 9766 8954 9818
rect 8966 9766 9018 9818
rect 9030 9766 9082 9818
rect 2964 9664 3016 9716
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 2964 9571 3016 9580
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 3424 9528 3476 9580
rect 3884 9596 3936 9648
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 4160 9528 4212 9580
rect 3884 9460 3936 9512
rect 4528 9528 4580 9580
rect 4068 9392 4120 9444
rect 4620 9392 4672 9444
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 6368 9528 6420 9580
rect 4988 9392 5040 9444
rect 3424 9324 3476 9376
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 5908 9392 5960 9444
rect 7748 9596 7800 9648
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 7472 9528 7524 9537
rect 7656 9460 7708 9512
rect 7840 9528 7892 9580
rect 8576 9460 8628 9512
rect 1973 9222 2025 9274
rect 2037 9222 2089 9274
rect 2101 9222 2153 9274
rect 2165 9222 2217 9274
rect 2229 9222 2281 9274
rect 4020 9222 4072 9274
rect 4084 9222 4136 9274
rect 4148 9222 4200 9274
rect 4212 9222 4264 9274
rect 4276 9222 4328 9274
rect 6067 9222 6119 9274
rect 6131 9222 6183 9274
rect 6195 9222 6247 9274
rect 6259 9222 6311 9274
rect 6323 9222 6375 9274
rect 8114 9222 8166 9274
rect 8178 9222 8230 9274
rect 8242 9222 8294 9274
rect 8306 9222 8358 9274
rect 8370 9222 8422 9274
rect 2872 9120 2924 9172
rect 4620 9120 4672 9172
rect 4896 9120 4948 9172
rect 5908 9120 5960 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 5724 8984 5776 9036
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 4528 8848 4580 8900
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 3148 8823 3200 8832
rect 3148 8789 3157 8823
rect 3157 8789 3191 8823
rect 3191 8789 3200 8823
rect 3148 8780 3200 8789
rect 5172 8780 5224 8832
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 7472 9052 7524 9104
rect 8576 9052 8628 9104
rect 6460 8916 6512 8968
rect 7104 8916 7156 8968
rect 7288 8916 7340 8968
rect 7380 8891 7432 8900
rect 7380 8857 7389 8891
rect 7389 8857 7423 8891
rect 7423 8857 7432 8891
rect 7380 8848 7432 8857
rect 2633 8678 2685 8730
rect 2697 8678 2749 8730
rect 2761 8678 2813 8730
rect 2825 8678 2877 8730
rect 2889 8678 2941 8730
rect 4680 8678 4732 8730
rect 4744 8678 4796 8730
rect 4808 8678 4860 8730
rect 4872 8678 4924 8730
rect 4936 8678 4988 8730
rect 6727 8678 6779 8730
rect 6791 8678 6843 8730
rect 6855 8678 6907 8730
rect 6919 8678 6971 8730
rect 6983 8678 7035 8730
rect 8774 8678 8826 8730
rect 8838 8678 8890 8730
rect 8902 8678 8954 8730
rect 8966 8678 9018 8730
rect 9030 8678 9082 8730
rect 8484 8576 8536 8628
rect 5172 8508 5224 8560
rect 7104 8508 7156 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 6920 8440 6972 8492
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 3240 8236 3292 8288
rect 1973 8134 2025 8186
rect 2037 8134 2089 8186
rect 2101 8134 2153 8186
rect 2165 8134 2217 8186
rect 2229 8134 2281 8186
rect 4020 8134 4072 8186
rect 4084 8134 4136 8186
rect 4148 8134 4200 8186
rect 4212 8134 4264 8186
rect 4276 8134 4328 8186
rect 6067 8134 6119 8186
rect 6131 8134 6183 8186
rect 6195 8134 6247 8186
rect 6259 8134 6311 8186
rect 6323 8134 6375 8186
rect 8114 8134 8166 8186
rect 8178 8134 8230 8186
rect 8242 8134 8294 8186
rect 8306 8134 8358 8186
rect 8370 8134 8422 8186
rect 3240 8032 3292 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 6920 8032 6972 8084
rect 3056 7964 3108 8016
rect 3240 7828 3292 7880
rect 3516 7896 3568 7948
rect 7472 7896 7524 7948
rect 1400 7735 1452 7744
rect 1400 7701 1409 7735
rect 1409 7701 1443 7735
rect 1443 7701 1452 7735
rect 1400 7692 1452 7701
rect 2964 7692 3016 7744
rect 3608 7692 3660 7744
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 3792 7803 3844 7812
rect 3792 7769 3801 7803
rect 3801 7769 3835 7803
rect 3835 7769 3844 7803
rect 3792 7760 3844 7769
rect 3884 7760 3936 7812
rect 9220 7828 9272 7880
rect 5724 7760 5776 7812
rect 8484 7803 8536 7812
rect 8484 7769 8493 7803
rect 8493 7769 8527 7803
rect 8527 7769 8536 7803
rect 8484 7760 8536 7769
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5264 7692 5316 7701
rect 5448 7692 5500 7744
rect 2633 7590 2685 7642
rect 2697 7590 2749 7642
rect 2761 7590 2813 7642
rect 2825 7590 2877 7642
rect 2889 7590 2941 7642
rect 4680 7590 4732 7642
rect 4744 7590 4796 7642
rect 4808 7590 4860 7642
rect 4872 7590 4924 7642
rect 4936 7590 4988 7642
rect 6727 7590 6779 7642
rect 6791 7590 6843 7642
rect 6855 7590 6907 7642
rect 6919 7590 6971 7642
rect 6983 7590 7035 7642
rect 8774 7590 8826 7642
rect 8838 7590 8890 7642
rect 8902 7590 8954 7642
rect 8966 7590 9018 7642
rect 9030 7590 9082 7642
rect 2964 7488 3016 7540
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 5264 7488 5316 7540
rect 1584 7420 1636 7472
rect 2412 7420 2464 7472
rect 3332 7352 3384 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 5816 7488 5868 7540
rect 6644 7420 6696 7472
rect 4436 7284 4488 7336
rect 5264 7284 5316 7336
rect 4620 7216 4672 7268
rect 5632 7216 5684 7268
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 8024 7420 8076 7472
rect 8668 7420 8720 7472
rect 2320 7148 2372 7200
rect 5816 7148 5868 7200
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 7932 7148 7984 7200
rect 1973 7046 2025 7098
rect 2037 7046 2089 7098
rect 2101 7046 2153 7098
rect 2165 7046 2217 7098
rect 2229 7046 2281 7098
rect 4020 7046 4072 7098
rect 4084 7046 4136 7098
rect 4148 7046 4200 7098
rect 4212 7046 4264 7098
rect 4276 7046 4328 7098
rect 6067 7046 6119 7098
rect 6131 7046 6183 7098
rect 6195 7046 6247 7098
rect 6259 7046 6311 7098
rect 6323 7046 6375 7098
rect 8114 7046 8166 7098
rect 8178 7046 8230 7098
rect 8242 7046 8294 7098
rect 8306 7046 8358 7098
rect 8370 7046 8422 7098
rect 3240 6987 3292 6996
rect 3240 6953 3249 6987
rect 3249 6953 3283 6987
rect 3283 6953 3292 6987
rect 3240 6944 3292 6953
rect 3792 6944 3844 6996
rect 5448 6944 5500 6996
rect 5540 6987 5592 6996
rect 5540 6953 5549 6987
rect 5549 6953 5583 6987
rect 5583 6953 5592 6987
rect 5540 6944 5592 6953
rect 5724 6944 5776 6996
rect 6000 6944 6052 6996
rect 7840 6944 7892 6996
rect 1584 6808 1636 6860
rect 3148 6808 3200 6860
rect 5908 6876 5960 6928
rect 4620 6808 4672 6860
rect 7932 6876 7984 6928
rect 3056 6740 3108 6792
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 3240 6715 3292 6724
rect 3240 6681 3249 6715
rect 3249 6681 3283 6715
rect 3283 6681 3292 6715
rect 3240 6672 3292 6681
rect 3424 6672 3476 6724
rect 4436 6672 4488 6724
rect 5540 6715 5592 6724
rect 5540 6681 5549 6715
rect 5549 6681 5583 6715
rect 5583 6681 5592 6715
rect 5540 6672 5592 6681
rect 6644 6740 6696 6792
rect 7656 6740 7708 6792
rect 8024 6808 8076 6860
rect 7564 6672 7616 6724
rect 7748 6672 7800 6724
rect 3608 6604 3660 6656
rect 3792 6604 3844 6656
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 5080 6604 5132 6656
rect 5816 6604 5868 6656
rect 7104 6604 7156 6656
rect 7288 6604 7340 6656
rect 8668 6740 8720 6792
rect 8576 6604 8628 6656
rect 2633 6502 2685 6554
rect 2697 6502 2749 6554
rect 2761 6502 2813 6554
rect 2825 6502 2877 6554
rect 2889 6502 2941 6554
rect 4680 6502 4732 6554
rect 4744 6502 4796 6554
rect 4808 6502 4860 6554
rect 4872 6502 4924 6554
rect 4936 6502 4988 6554
rect 6727 6502 6779 6554
rect 6791 6502 6843 6554
rect 6855 6502 6907 6554
rect 6919 6502 6971 6554
rect 6983 6502 7035 6554
rect 8774 6502 8826 6554
rect 8838 6502 8890 6554
rect 8902 6502 8954 6554
rect 8966 6502 9018 6554
rect 9030 6502 9082 6554
rect 2320 6400 2372 6452
rect 3056 6400 3108 6452
rect 3240 6400 3292 6452
rect 2412 6332 2464 6384
rect 3424 6332 3476 6384
rect 5080 6332 5132 6384
rect 5172 6375 5224 6384
rect 5172 6341 5181 6375
rect 5181 6341 5215 6375
rect 5215 6341 5224 6375
rect 5172 6332 5224 6341
rect 1860 6264 1912 6316
rect 3884 6307 3936 6316
rect 2320 6171 2372 6180
rect 2320 6137 2329 6171
rect 2329 6137 2363 6171
rect 2363 6137 2372 6171
rect 2320 6128 2372 6137
rect 3884 6273 3888 6307
rect 3888 6273 3922 6307
rect 3922 6273 3936 6307
rect 3884 6264 3936 6273
rect 4252 6307 4304 6316
rect 3608 6196 3660 6248
rect 4252 6273 4260 6307
rect 4260 6273 4294 6307
rect 4294 6273 4304 6307
rect 4252 6264 4304 6273
rect 4528 6264 4580 6316
rect 7564 6400 7616 6452
rect 7288 6332 7340 6384
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 7472 6264 7524 6316
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 1584 6060 1636 6112
rect 1860 6060 1912 6112
rect 3056 6128 3108 6180
rect 5172 6128 5224 6180
rect 5724 6128 5776 6180
rect 6000 6128 6052 6180
rect 7932 6128 7984 6180
rect 5540 6060 5592 6112
rect 5816 6060 5868 6112
rect 7748 6060 7800 6112
rect 8024 6060 8076 6112
rect 1973 5958 2025 6010
rect 2037 5958 2089 6010
rect 2101 5958 2153 6010
rect 2165 5958 2217 6010
rect 2229 5958 2281 6010
rect 4020 5958 4072 6010
rect 4084 5958 4136 6010
rect 4148 5958 4200 6010
rect 4212 5958 4264 6010
rect 4276 5958 4328 6010
rect 6067 5958 6119 6010
rect 6131 5958 6183 6010
rect 6195 5958 6247 6010
rect 6259 5958 6311 6010
rect 6323 5958 6375 6010
rect 8114 5958 8166 6010
rect 8178 5958 8230 6010
rect 8242 5958 8294 6010
rect 8306 5958 8358 6010
rect 8370 5958 8422 6010
rect 4528 5856 4580 5908
rect 3516 5720 3568 5772
rect 5264 5788 5316 5840
rect 5908 5788 5960 5840
rect 6552 5831 6604 5840
rect 6552 5797 6561 5831
rect 6561 5797 6595 5831
rect 6595 5797 6604 5831
rect 6552 5788 6604 5797
rect 1400 5652 1452 5704
rect 2964 5652 3016 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4620 5652 4672 5704
rect 5540 5652 5592 5704
rect 7840 5831 7892 5840
rect 7840 5797 7849 5831
rect 7849 5797 7883 5831
rect 7883 5797 7892 5831
rect 7840 5788 7892 5797
rect 5264 5627 5316 5636
rect 5264 5593 5273 5627
rect 5273 5593 5307 5627
rect 5307 5593 5316 5627
rect 5264 5584 5316 5593
rect 6644 5516 6696 5568
rect 9312 5516 9364 5568
rect 2633 5414 2685 5466
rect 2697 5414 2749 5466
rect 2761 5414 2813 5466
rect 2825 5414 2877 5466
rect 2889 5414 2941 5466
rect 4680 5414 4732 5466
rect 4744 5414 4796 5466
rect 4808 5414 4860 5466
rect 4872 5414 4924 5466
rect 4936 5414 4988 5466
rect 6727 5414 6779 5466
rect 6791 5414 6843 5466
rect 6855 5414 6907 5466
rect 6919 5414 6971 5466
rect 6983 5414 7035 5466
rect 8774 5414 8826 5466
rect 8838 5414 8890 5466
rect 8902 5414 8954 5466
rect 8966 5414 9018 5466
rect 9030 5414 9082 5466
rect 2412 5312 2464 5364
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 3792 5312 3844 5364
rect 4160 5312 4212 5364
rect 4436 5312 4488 5364
rect 7564 5355 7616 5364
rect 7564 5321 7573 5355
rect 7573 5321 7607 5355
rect 7607 5321 7616 5355
rect 7564 5312 7616 5321
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3240 5219 3292 5228
rect 3240 5185 3248 5219
rect 3248 5185 3282 5219
rect 3282 5185 3292 5219
rect 3240 5176 3292 5185
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 4896 5176 4948 5228
rect 5080 5244 5132 5296
rect 5172 5287 5224 5296
rect 5172 5253 5181 5287
rect 5181 5253 5215 5287
rect 5215 5253 5224 5287
rect 5172 5244 5224 5253
rect 3884 5108 3936 5160
rect 5448 5176 5500 5228
rect 5540 5176 5592 5228
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 6644 5176 6696 5228
rect 7288 5176 7340 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 7656 5108 7708 5160
rect 2320 4972 2372 5024
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 1973 4870 2025 4922
rect 2037 4870 2089 4922
rect 2101 4870 2153 4922
rect 2165 4870 2217 4922
rect 2229 4870 2281 4922
rect 4020 4870 4072 4922
rect 4084 4870 4136 4922
rect 4148 4870 4200 4922
rect 4212 4870 4264 4922
rect 4276 4870 4328 4922
rect 6067 4870 6119 4922
rect 6131 4870 6183 4922
rect 6195 4870 6247 4922
rect 6259 4870 6311 4922
rect 6323 4870 6375 4922
rect 8114 4870 8166 4922
rect 8178 4870 8230 4922
rect 8242 4870 8294 4922
rect 8306 4870 8358 4922
rect 8370 4870 8422 4922
rect 3332 4768 3384 4820
rect 5356 4768 5408 4820
rect 6460 4768 6512 4820
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 5632 4700 5684 4752
rect 4528 4632 4580 4684
rect 3240 4496 3292 4548
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 7472 4564 7524 4616
rect 8668 4496 8720 4548
rect 5172 4428 5224 4480
rect 5448 4428 5500 4480
rect 2633 4326 2685 4378
rect 2697 4326 2749 4378
rect 2761 4326 2813 4378
rect 2825 4326 2877 4378
rect 2889 4326 2941 4378
rect 4680 4326 4732 4378
rect 4744 4326 4796 4378
rect 4808 4326 4860 4378
rect 4872 4326 4924 4378
rect 4936 4326 4988 4378
rect 6727 4326 6779 4378
rect 6791 4326 6843 4378
rect 6855 4326 6907 4378
rect 6919 4326 6971 4378
rect 6983 4326 7035 4378
rect 8774 4326 8826 4378
rect 8838 4326 8890 4378
rect 8902 4326 8954 4378
rect 8966 4326 9018 4378
rect 9030 4326 9082 4378
rect 5816 4224 5868 4276
rect 6644 4224 6696 4276
rect 4436 4156 4488 4208
rect 3884 4088 3936 4140
rect 6460 4156 6512 4208
rect 6368 4088 6420 4140
rect 3976 3952 4028 4004
rect 5172 3952 5224 4004
rect 8484 4088 8536 4140
rect 5908 3884 5960 3936
rect 6460 3884 6512 3936
rect 7288 4020 7340 4072
rect 1973 3782 2025 3834
rect 2037 3782 2089 3834
rect 2101 3782 2153 3834
rect 2165 3782 2217 3834
rect 2229 3782 2281 3834
rect 4020 3782 4072 3834
rect 4084 3782 4136 3834
rect 4148 3782 4200 3834
rect 4212 3782 4264 3834
rect 4276 3782 4328 3834
rect 6067 3782 6119 3834
rect 6131 3782 6183 3834
rect 6195 3782 6247 3834
rect 6259 3782 6311 3834
rect 6323 3782 6375 3834
rect 8114 3782 8166 3834
rect 8178 3782 8230 3834
rect 8242 3782 8294 3834
rect 8306 3782 8358 3834
rect 8370 3782 8422 3834
rect 1860 3680 1912 3732
rect 2320 3612 2372 3664
rect 3700 3680 3752 3732
rect 1492 3451 1544 3460
rect 1492 3417 1501 3451
rect 1501 3417 1535 3451
rect 1535 3417 1544 3451
rect 1492 3408 1544 3417
rect 940 3340 992 3392
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 5356 3476 5408 3528
rect 5540 3680 5592 3732
rect 5908 3680 5960 3732
rect 6552 3476 6604 3528
rect 5632 3408 5684 3460
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 5908 3340 5960 3392
rect 2633 3238 2685 3290
rect 2697 3238 2749 3290
rect 2761 3238 2813 3290
rect 2825 3238 2877 3290
rect 2889 3238 2941 3290
rect 4680 3238 4732 3290
rect 4744 3238 4796 3290
rect 4808 3238 4860 3290
rect 4872 3238 4924 3290
rect 4936 3238 4988 3290
rect 6727 3238 6779 3290
rect 6791 3238 6843 3290
rect 6855 3238 6907 3290
rect 6919 3238 6971 3290
rect 6983 3238 7035 3290
rect 8774 3238 8826 3290
rect 8838 3238 8890 3290
rect 8902 3238 8954 3290
rect 8966 3238 9018 3290
rect 9030 3238 9082 3290
rect 4528 3136 4580 3188
rect 5080 3136 5132 3188
rect 6460 3136 6512 3188
rect 6644 3136 6696 3188
rect 3700 3068 3752 3120
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 20 3000 72 3052
rect 5724 3000 5776 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 3056 2907 3108 2916
rect 3056 2873 3065 2907
rect 3065 2873 3099 2907
rect 3099 2873 3108 2907
rect 3056 2864 3108 2873
rect 4436 2839 4488 2848
rect 4436 2805 4445 2839
rect 4445 2805 4479 2839
rect 4479 2805 4488 2839
rect 4436 2796 4488 2805
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 8852 2839 8904 2848
rect 8852 2805 8861 2839
rect 8861 2805 8895 2839
rect 8895 2805 8904 2839
rect 8852 2796 8904 2805
rect 1973 2694 2025 2746
rect 2037 2694 2089 2746
rect 2101 2694 2153 2746
rect 2165 2694 2217 2746
rect 2229 2694 2281 2746
rect 4020 2694 4072 2746
rect 4084 2694 4136 2746
rect 4148 2694 4200 2746
rect 4212 2694 4264 2746
rect 4276 2694 4328 2746
rect 6067 2694 6119 2746
rect 6131 2694 6183 2746
rect 6195 2694 6247 2746
rect 6259 2694 6311 2746
rect 6323 2694 6375 2746
rect 8114 2694 8166 2746
rect 8178 2694 8230 2746
rect 8242 2694 8294 2746
rect 8306 2694 8358 2746
rect 8370 2694 8422 2746
rect 1492 2592 1544 2644
rect 4436 2592 4488 2644
rect 3056 2456 3108 2508
rect 5632 2592 5684 2644
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 8668 2592 8720 2644
rect 3424 2388 3476 2440
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 7748 2388 7800 2440
rect 10324 2388 10376 2440
rect 3516 2252 3568 2304
rect 2633 2150 2685 2202
rect 2697 2150 2749 2202
rect 2761 2150 2813 2202
rect 2825 2150 2877 2202
rect 2889 2150 2941 2202
rect 4680 2150 4732 2202
rect 4744 2150 4796 2202
rect 4808 2150 4860 2202
rect 4872 2150 4924 2202
rect 4936 2150 4988 2202
rect 6727 2150 6779 2202
rect 6791 2150 6843 2202
rect 6855 2150 6907 2202
rect 6919 2150 6971 2202
rect 6983 2150 7035 2202
rect 8774 2150 8826 2202
rect 8838 2150 8890 2202
rect 8902 2150 8954 2202
rect 8966 2150 9018 2202
rect 9030 2150 9082 2202
<< metal2 >>
rect 1306 11817 1362 12617
rect 3882 11817 3938 12617
rect 6458 11817 6514 12617
rect 9034 11817 9090 12617
rect 938 10976 994 10985
rect 938 10911 994 10920
rect 952 10062 980 10911
rect 1320 10266 1348 11817
rect 1973 10364 2281 10373
rect 1973 10362 1979 10364
rect 2035 10362 2059 10364
rect 2115 10362 2139 10364
rect 2195 10362 2219 10364
rect 2275 10362 2281 10364
rect 2035 10310 2037 10362
rect 2217 10310 2219 10362
rect 1973 10308 1979 10310
rect 2035 10308 2059 10310
rect 2115 10308 2139 10310
rect 2195 10308 2219 10310
rect 2275 10308 2281 10310
rect 1973 10299 2281 10308
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 940 10056 992 10062
rect 940 9998 992 10004
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1584 8288 1636 8294
rect 1398 8256 1454 8265
rect 1584 8230 1636 8236
rect 1398 8191 1454 8200
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1412 5710 1440 7686
rect 1596 7478 1624 8230
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1596 6866 1624 7414
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6118 1624 6802
rect 1872 6322 1900 9862
rect 2633 9820 2941 9829
rect 2633 9818 2639 9820
rect 2695 9818 2719 9820
rect 2775 9818 2799 9820
rect 2855 9818 2879 9820
rect 2935 9818 2941 9820
rect 2695 9766 2697 9818
rect 2877 9766 2879 9818
rect 2633 9764 2639 9766
rect 2695 9764 2719 9766
rect 2775 9764 2799 9766
rect 2855 9764 2879 9766
rect 2935 9764 2941 9766
rect 2633 9755 2941 9764
rect 2976 9722 3004 10134
rect 3896 10062 3924 11817
rect 4020 10364 4328 10373
rect 4020 10362 4026 10364
rect 4082 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4328 10364
rect 4082 10310 4084 10362
rect 4264 10310 4266 10362
rect 4020 10308 4026 10310
rect 4082 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4328 10310
rect 4020 10299 4328 10308
rect 6067 10364 6375 10373
rect 6067 10362 6073 10364
rect 6129 10362 6153 10364
rect 6209 10362 6233 10364
rect 6289 10362 6313 10364
rect 6369 10362 6375 10364
rect 6129 10310 6131 10362
rect 6311 10310 6313 10362
rect 6067 10308 6073 10310
rect 6129 10308 6153 10310
rect 6209 10308 6233 10310
rect 6289 10308 6313 10310
rect 6369 10308 6375 10310
rect 6067 10299 6375 10308
rect 6472 10062 6500 11817
rect 8114 10364 8422 10373
rect 8114 10362 8120 10364
rect 8176 10362 8200 10364
rect 8256 10362 8280 10364
rect 8336 10362 8360 10364
rect 8416 10362 8422 10364
rect 8176 10310 8178 10362
rect 8358 10310 8360 10362
rect 8114 10308 8120 10310
rect 8176 10308 8200 10310
rect 8256 10308 8280 10310
rect 8336 10308 8360 10310
rect 8416 10308 8422 10310
rect 8114 10299 8422 10308
rect 9048 10266 9076 11817
rect 9218 10976 9274 10985
rect 9218 10911 9274 10920
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9232 10062 9260 10911
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 4680 9820 4988 9829
rect 4680 9818 4686 9820
rect 4742 9818 4766 9820
rect 4822 9818 4846 9820
rect 4902 9818 4926 9820
rect 4982 9818 4988 9820
rect 4742 9766 4744 9818
rect 4924 9766 4926 9818
rect 4680 9764 4686 9766
rect 4742 9764 4766 9766
rect 4822 9764 4846 9766
rect 4902 9764 4926 9766
rect 4982 9764 4988 9766
rect 4680 9755 4988 9764
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 2976 9586 3004 9658
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3436 9382 3464 9522
rect 3896 9518 3924 9590
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 1973 9276 2281 9285
rect 1973 9274 1979 9276
rect 2035 9274 2059 9276
rect 2115 9274 2139 9276
rect 2195 9274 2219 9276
rect 2275 9274 2281 9276
rect 2035 9222 2037 9274
rect 2217 9222 2219 9274
rect 1973 9220 1979 9222
rect 2035 9220 2059 9222
rect 2115 9220 2139 9222
rect 2195 9220 2219 9222
rect 2275 9220 2281 9222
rect 1973 9211 2281 9220
rect 2884 9178 2912 9318
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 2633 8732 2941 8741
rect 2633 8730 2639 8732
rect 2695 8730 2719 8732
rect 2775 8730 2799 8732
rect 2855 8730 2879 8732
rect 2935 8730 2941 8732
rect 2695 8678 2697 8730
rect 2877 8678 2879 8730
rect 2633 8676 2639 8678
rect 2695 8676 2719 8678
rect 2775 8676 2799 8678
rect 2855 8676 2879 8678
rect 2935 8676 2941 8678
rect 2633 8667 2941 8676
rect 1973 8188 2281 8197
rect 1973 8186 1979 8188
rect 2035 8186 2059 8188
rect 2115 8186 2139 8188
rect 2195 8186 2219 8188
rect 2275 8186 2281 8188
rect 2035 8134 2037 8186
rect 2217 8134 2219 8186
rect 1973 8132 1979 8134
rect 2035 8132 2059 8134
rect 2115 8132 2139 8134
rect 2195 8132 2219 8134
rect 2275 8132 2281 8134
rect 1973 8123 2281 8132
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2633 7644 2941 7653
rect 2633 7642 2639 7644
rect 2695 7642 2719 7644
rect 2775 7642 2799 7644
rect 2855 7642 2879 7644
rect 2935 7642 2941 7644
rect 2695 7590 2697 7642
rect 2877 7590 2879 7642
rect 2633 7588 2639 7590
rect 2695 7588 2719 7590
rect 2775 7588 2799 7590
rect 2855 7588 2879 7590
rect 2935 7588 2941 7590
rect 2633 7579 2941 7588
rect 2976 7546 3004 7686
rect 3068 7546 3096 7958
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 1973 7100 2281 7109
rect 1973 7098 1979 7100
rect 2035 7098 2059 7100
rect 2115 7098 2139 7100
rect 2195 7098 2219 7100
rect 2275 7098 2281 7100
rect 2035 7046 2037 7098
rect 2217 7046 2219 7098
rect 1973 7044 1979 7046
rect 2035 7044 2059 7046
rect 2115 7044 2139 7046
rect 2195 7044 2219 7046
rect 2275 7044 2281 7046
rect 1973 7035 2281 7044
rect 2332 6458 2360 7142
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 2332 6186 2360 6394
rect 2424 6390 2452 7414
rect 3160 6866 3188 8774
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 8090 3280 8230
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7002 3280 7822
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2633 6556 2941 6565
rect 2633 6554 2639 6556
rect 2695 6554 2719 6556
rect 2775 6554 2799 6556
rect 2855 6554 2879 6556
rect 2935 6554 2941 6556
rect 2695 6502 2697 6554
rect 2877 6502 2879 6554
rect 2633 6500 2639 6502
rect 2695 6500 2719 6502
rect 2775 6500 2799 6502
rect 2855 6500 2879 6502
rect 2935 6500 2941 6502
rect 2633 6491 2941 6500
rect 3068 6458 3096 6734
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3252 6458 3280 6666
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 2412 6384 2464 6390
rect 3344 6338 3372 7346
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3436 6390 3464 6666
rect 2412 6326 2464 6332
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1582 5471 1638 5480
rect 1872 5234 1900 6054
rect 1973 6012 2281 6021
rect 1973 6010 1979 6012
rect 2035 6010 2059 6012
rect 2115 6010 2139 6012
rect 2195 6010 2219 6012
rect 2275 6010 2281 6012
rect 2035 5958 2037 6010
rect 2217 5958 2219 6010
rect 1973 5956 1979 5958
rect 2035 5956 2059 5958
rect 2115 5956 2139 5958
rect 2195 5956 2219 5958
rect 2275 5956 2281 5958
rect 1973 5947 2281 5956
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1872 3738 1900 5170
rect 2332 5030 2360 6122
rect 2424 5370 2452 6326
rect 3252 6310 3372 6338
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2633 5468 2941 5477
rect 2633 5466 2639 5468
rect 2695 5466 2719 5468
rect 2775 5466 2799 5468
rect 2855 5466 2879 5468
rect 2935 5466 2941 5468
rect 2695 5414 2697 5466
rect 2877 5414 2879 5466
rect 2633 5412 2639 5414
rect 2695 5412 2719 5414
rect 2775 5412 2799 5414
rect 2855 5412 2879 5414
rect 2935 5412 2941 5414
rect 2633 5403 2941 5412
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2976 5234 3004 5646
rect 3068 5234 3096 6122
rect 3252 5234 3280 6310
rect 3528 5778 3556 7890
rect 3896 7818 3924 9454
rect 4068 9444 4120 9450
rect 4172 9432 4200 9522
rect 4120 9404 4200 9432
rect 4068 9386 4120 9392
rect 4020 9276 4328 9285
rect 4020 9274 4026 9276
rect 4082 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4328 9276
rect 4082 9222 4084 9274
rect 4264 9222 4266 9274
rect 4020 9220 4026 9222
rect 4082 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4328 9222
rect 4020 9211 4328 9220
rect 4540 8906 4568 9522
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4632 9178 4660 9386
rect 4908 9178 4936 9658
rect 5632 9580 5684 9586
rect 6000 9580 6052 9586
rect 5632 9522 5684 9528
rect 5828 9540 6000 9568
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5000 8974 5028 9386
rect 5644 8974 5672 9522
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 9042 5764 9318
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4680 8732 4988 8741
rect 4680 8730 4686 8732
rect 4742 8730 4766 8732
rect 4822 8730 4846 8732
rect 4902 8730 4926 8732
rect 4982 8730 4988 8732
rect 4742 8678 4744 8730
rect 4924 8678 4926 8730
rect 4680 8676 4686 8678
rect 4742 8676 4766 8678
rect 4822 8676 4846 8678
rect 4902 8676 4926 8678
rect 4982 8676 4988 8678
rect 4680 8667 4988 8676
rect 5184 8566 5212 8774
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 4020 8188 4328 8197
rect 4020 8186 4026 8188
rect 4082 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4328 8188
rect 4082 8134 4084 8186
rect 4264 8134 4266 8186
rect 4020 8132 4026 8134
rect 4082 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4328 8134
rect 4020 8123 4328 8132
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3608 7744 3660 7750
rect 3804 7698 3832 7754
rect 3660 7692 3832 7698
rect 3608 7686 3832 7692
rect 3620 7670 3832 7686
rect 3804 7018 3832 7670
rect 3712 7002 3832 7018
rect 3712 6996 3844 7002
rect 3712 6990 3792 6996
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6254 3648 6598
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3620 5370 3648 6190
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1973 4924 2281 4933
rect 1973 4922 1979 4924
rect 2035 4922 2059 4924
rect 2115 4922 2139 4924
rect 2195 4922 2219 4924
rect 2275 4922 2281 4924
rect 2035 4870 2037 4922
rect 2217 4870 2219 4922
rect 1973 4868 1979 4870
rect 2035 4868 2059 4870
rect 2115 4868 2139 4870
rect 2195 4868 2219 4870
rect 2275 4868 2281 4870
rect 1973 4859 2281 4868
rect 1973 3836 2281 3845
rect 1973 3834 1979 3836
rect 2035 3834 2059 3836
rect 2115 3834 2139 3836
rect 2195 3834 2219 3836
rect 2275 3834 2281 3836
rect 2035 3782 2037 3834
rect 2217 3782 2219 3834
rect 1973 3780 1979 3782
rect 2035 3780 2059 3782
rect 2115 3780 2139 3782
rect 2195 3780 2219 3782
rect 2275 3780 2281 3782
rect 1973 3771 2281 3780
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2332 3670 2360 4966
rect 3252 4554 3280 5170
rect 3344 4826 3372 5170
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 2633 4380 2941 4389
rect 2633 4378 2639 4380
rect 2695 4378 2719 4380
rect 2775 4378 2799 4380
rect 2855 4378 2879 4380
rect 2935 4378 2941 4380
rect 2695 4326 2697 4378
rect 2877 4326 2879 4378
rect 2633 4324 2639 4326
rect 2695 4324 2719 4326
rect 2775 4324 2799 4326
rect 2855 4324 2879 4326
rect 2935 4324 2941 4326
rect 2633 4315 2941 4324
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 940 3392 992 3398
rect 940 3334 992 3340
rect 20 3052 72 3058
rect 20 2994 72 3000
rect 32 800 60 2994
rect 952 2825 980 3334
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 1504 2650 1532 3402
rect 2633 3292 2941 3301
rect 2633 3290 2639 3292
rect 2695 3290 2719 3292
rect 2775 3290 2799 3292
rect 2855 3290 2879 3292
rect 2935 3290 2941 3292
rect 2695 3238 2697 3290
rect 2877 3238 2879 3290
rect 2633 3236 2639 3238
rect 2695 3236 2719 3238
rect 2775 3236 2799 3238
rect 2855 3236 2879 3238
rect 2935 3236 2941 3238
rect 2633 3227 2941 3236
rect 2502 2952 2558 2961
rect 2502 2887 2558 2896
rect 3056 2916 3108 2922
rect 1973 2748 2281 2757
rect 1973 2746 1979 2748
rect 2035 2746 2059 2748
rect 2115 2746 2139 2748
rect 2195 2746 2219 2748
rect 2275 2746 2281 2748
rect 2035 2694 2037 2746
rect 2217 2694 2219 2746
rect 1973 2692 1979 2694
rect 2035 2692 2059 2694
rect 2115 2692 2139 2694
rect 2195 2692 2219 2694
rect 2275 2692 2281 2694
rect 1973 2683 2281 2692
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 2516 1986 2544 2887
rect 3056 2858 3108 2864
rect 3068 2514 3096 2858
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3436 2446 3464 4966
rect 3712 3738 3740 6990
rect 3792 6938 3844 6944
rect 3792 6656 3844 6662
rect 3896 6644 3924 7754
rect 4680 7644 4988 7653
rect 4680 7642 4686 7644
rect 4742 7642 4766 7644
rect 4822 7642 4846 7644
rect 4902 7642 4926 7644
rect 4982 7642 4988 7644
rect 4742 7590 4744 7642
rect 4924 7590 4926 7642
rect 4680 7588 4686 7590
rect 4742 7588 4766 7590
rect 4822 7588 4846 7590
rect 4902 7588 4926 7590
rect 4982 7588 4988 7590
rect 4680 7579 4988 7588
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4020 7100 4328 7109
rect 4020 7098 4026 7100
rect 4082 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4328 7100
rect 4082 7046 4084 7098
rect 4264 7046 4266 7098
rect 4020 7044 4026 7046
rect 4082 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4328 7046
rect 4020 7035 4328 7044
rect 3844 6616 3924 6644
rect 4252 6656 4304 6662
rect 3792 6598 3844 6604
rect 4252 6598 4304 6604
rect 3804 5710 3832 6598
rect 4264 6322 4292 6598
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3804 4604 3832 5306
rect 3896 5166 3924 6258
rect 4020 6012 4328 6021
rect 4020 6010 4026 6012
rect 4082 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4328 6012
rect 4082 5958 4084 6010
rect 4264 5958 4266 6010
rect 4020 5956 4026 5958
rect 4082 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4328 5958
rect 4020 5947 4328 5956
rect 4158 5808 4214 5817
rect 4158 5743 4214 5752
rect 4172 5710 4200 5743
rect 4160 5704 4212 5710
rect 4356 5681 4384 7346
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4448 6730 4476 7278
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4632 6866 4660 7210
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4680 6556 4988 6565
rect 4680 6554 4686 6556
rect 4742 6554 4766 6556
rect 4822 6554 4846 6556
rect 4902 6554 4926 6556
rect 4982 6554 4988 6556
rect 4742 6502 4744 6554
rect 4924 6502 4926 6554
rect 4680 6500 4686 6502
rect 4742 6500 4766 6502
rect 4822 6500 4846 6502
rect 4902 6500 4926 6502
rect 4982 6500 4988 6502
rect 4680 6491 4988 6500
rect 5092 6390 5120 6598
rect 5184 6390 5212 7822
rect 5460 7750 5488 8774
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5276 7546 5304 7686
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4540 5914 4568 6258
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4620 5704 4672 5710
rect 4160 5646 4212 5652
rect 4342 5672 4398 5681
rect 4172 5370 4200 5646
rect 4342 5607 4398 5616
rect 4448 5664 4620 5692
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 4020 4924 4328 4933
rect 4020 4922 4026 4924
rect 4082 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4328 4924
rect 4082 4870 4084 4922
rect 4264 4870 4266 4922
rect 4020 4868 4026 4870
rect 4082 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4328 4870
rect 4020 4859 4328 4868
rect 3976 4616 4028 4622
rect 3804 4576 3976 4604
rect 3976 4558 4028 4564
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3700 3732 3752 3738
rect 3896 3720 3924 4082
rect 3988 4010 4016 4558
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 4020 3836 4328 3845
rect 4020 3834 4026 3836
rect 4082 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4328 3836
rect 4082 3782 4084 3834
rect 4264 3782 4266 3834
rect 4020 3780 4026 3782
rect 4082 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4328 3782
rect 4020 3771 4328 3780
rect 3896 3692 4200 3720
rect 3700 3674 3752 3680
rect 3712 3126 3740 3674
rect 4172 3534 4200 3692
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3712 2774 3740 3062
rect 3528 2746 3740 2774
rect 3804 2774 3832 3334
rect 4356 3126 4384 5607
rect 4448 5370 4476 5664
rect 4620 5646 4672 5652
rect 4680 5468 4988 5477
rect 4680 5466 4686 5468
rect 4742 5466 4766 5468
rect 4822 5466 4846 5468
rect 4902 5466 4926 5468
rect 4982 5466 4988 5468
rect 4742 5414 4744 5466
rect 4924 5414 4926 5466
rect 4680 5412 4686 5414
rect 4742 5412 4766 5414
rect 4822 5412 4846 5414
rect 4902 5412 4926 5414
rect 4982 5412 4988 5414
rect 4680 5403 4988 5412
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4448 4622 4476 5306
rect 5184 5302 5212 6122
rect 5276 5846 5304 7278
rect 5552 7002 5580 8026
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5460 6882 5488 6938
rect 5460 6854 5580 6882
rect 5552 6730 5580 6854
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5264 5840 5316 5846
rect 5316 5800 5396 5828
rect 5460 5817 5488 6258
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5264 5782 5316 5788
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5080 5296 5132 5302
rect 4894 5264 4950 5273
rect 5080 5238 5132 5244
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 4894 5199 4896 5208
rect 4948 5199 4950 5208
rect 4896 5170 4948 5176
rect 5092 4706 5120 5238
rect 5170 4720 5226 4729
rect 4528 4684 4580 4690
rect 5092 4678 5170 4706
rect 5170 4655 5226 4664
rect 4528 4626 4580 4632
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4448 4214 4476 4558
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4540 3194 4568 4626
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4680 4380 4988 4389
rect 4680 4378 4686 4380
rect 4742 4378 4766 4380
rect 4822 4378 4846 4380
rect 4902 4378 4926 4380
rect 4982 4378 4988 4380
rect 4742 4326 4744 4378
rect 4924 4326 4926 4378
rect 4680 4324 4686 4326
rect 4742 4324 4766 4326
rect 4822 4324 4846 4326
rect 4902 4324 4926 4326
rect 4982 4324 4988 4326
rect 4680 4315 4988 4324
rect 5184 4128 5212 4422
rect 5092 4100 5212 4128
rect 4680 3292 4988 3301
rect 4680 3290 4686 3292
rect 4742 3290 4766 3292
rect 4822 3290 4846 3292
rect 4902 3290 4926 3292
rect 4982 3290 4988 3292
rect 4742 3238 4744 3290
rect 4924 3238 4926 3290
rect 4680 3236 4686 3238
rect 4742 3236 4766 3238
rect 4822 3236 4846 3238
rect 4902 3236 4926 3238
rect 4982 3236 4988 3238
rect 4680 3227 4988 3236
rect 5092 3194 5120 4100
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5184 3398 5212 3946
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 5276 2961 5304 5578
rect 5368 4826 5396 5800
rect 5446 5808 5502 5817
rect 5446 5743 5502 5752
rect 5552 5710 5580 6054
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5234 5580 5646
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5368 3534 5396 4762
rect 5460 4486 5488 5170
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5552 3738 5580 4966
rect 5644 4758 5672 7210
rect 5736 7002 5764 7754
rect 5828 7546 5856 9540
rect 6368 9580 6420 9586
rect 6052 9540 6368 9568
rect 6000 9522 6052 9528
rect 6368 9522 6420 9528
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5920 9178 5948 9386
rect 6067 9276 6375 9285
rect 6067 9274 6073 9276
rect 6129 9274 6153 9276
rect 6209 9274 6233 9276
rect 6289 9274 6313 9276
rect 6369 9274 6375 9276
rect 6129 9222 6131 9274
rect 6311 9222 6313 9274
rect 6067 9220 6073 9222
rect 6129 9220 6153 9222
rect 6209 9220 6233 9222
rect 6289 9220 6313 9222
rect 6369 9220 6375 9222
rect 6067 9211 6375 9220
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6067 8188 6375 8197
rect 6067 8186 6073 8188
rect 6129 8186 6153 8188
rect 6209 8186 6233 8188
rect 6289 8186 6313 8188
rect 6369 8186 6375 8188
rect 6129 8134 6131 8186
rect 6311 8134 6313 8186
rect 6067 8132 6073 8134
rect 6129 8132 6153 8134
rect 6209 8132 6233 8134
rect 6289 8132 6313 8134
rect 6369 8132 6375 8134
rect 6067 8123 6375 8132
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6322 5764 6734
rect 5828 6662 5856 7142
rect 5920 6934 5948 7346
rect 6067 7100 6375 7109
rect 6067 7098 6073 7100
rect 6129 7098 6153 7100
rect 6209 7098 6233 7100
rect 6289 7098 6313 7100
rect 6369 7098 6375 7100
rect 6129 7046 6131 7098
rect 6311 7046 6313 7098
rect 6067 7044 6073 7046
rect 6129 7044 6153 7046
rect 6209 7044 6233 7046
rect 6289 7044 6313 7046
rect 6369 7044 6375 7046
rect 6067 7035 6375 7044
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5644 3466 5672 4694
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5736 3058 5764 6122
rect 5828 6118 5856 6598
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5920 5846 5948 6870
rect 6012 6186 6040 6938
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6067 6012 6375 6021
rect 6067 6010 6073 6012
rect 6129 6010 6153 6012
rect 6209 6010 6233 6012
rect 6289 6010 6313 6012
rect 6369 6010 6375 6012
rect 6129 5958 6131 6010
rect 6311 5958 6313 6010
rect 6067 5956 6073 5958
rect 6129 5956 6153 5958
rect 6209 5956 6233 5958
rect 6289 5956 6313 5958
rect 6369 5956 6375 5958
rect 6067 5947 6375 5956
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5920 5234 5948 5782
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6067 4924 6375 4933
rect 6067 4922 6073 4924
rect 6129 4922 6153 4924
rect 6209 4922 6233 4924
rect 6289 4922 6313 4924
rect 6369 4922 6375 4924
rect 6129 4870 6131 4922
rect 6311 4870 6313 4922
rect 6067 4868 6073 4870
rect 6129 4868 6153 4870
rect 6209 4868 6233 4870
rect 6289 4868 6313 4870
rect 6369 4868 6375 4870
rect 6067 4859 6375 4868
rect 6472 4826 6500 8910
rect 6656 7478 6684 9862
rect 6727 9820 7035 9829
rect 6727 9818 6733 9820
rect 6789 9818 6813 9820
rect 6869 9818 6893 9820
rect 6949 9818 6973 9820
rect 7029 9818 7035 9820
rect 6789 9766 6791 9818
rect 6971 9766 6973 9818
rect 6727 9764 6733 9766
rect 6789 9764 6813 9766
rect 6869 9764 6893 9766
rect 6949 9764 6973 9766
rect 7029 9764 7035 9766
rect 6727 9755 7035 9764
rect 7116 8974 7144 9930
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7484 9110 7512 9522
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7668 9058 7696 9454
rect 7760 9178 7788 9590
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7852 9058 7880 9522
rect 8114 9276 8422 9285
rect 8114 9274 8120 9276
rect 8176 9274 8200 9276
rect 8256 9274 8280 9276
rect 8336 9274 8360 9276
rect 8416 9274 8422 9276
rect 8176 9222 8178 9274
rect 8358 9222 8360 9274
rect 8114 9220 8120 9222
rect 8176 9220 8200 9222
rect 8256 9220 8280 9222
rect 8336 9220 8360 9222
rect 8416 9220 8422 9222
rect 8114 9211 8422 9220
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 6727 8732 7035 8741
rect 6727 8730 6733 8732
rect 6789 8730 6813 8732
rect 6869 8730 6893 8732
rect 6949 8730 6973 8732
rect 7029 8730 7035 8732
rect 6789 8678 6791 8730
rect 6971 8678 6973 8730
rect 6727 8676 6733 8678
rect 6789 8676 6813 8678
rect 6869 8676 6893 8678
rect 6949 8676 6973 8678
rect 7029 8676 7035 8678
rect 6727 8667 7035 8676
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6932 8090 6960 8434
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6727 7644 7035 7653
rect 6727 7642 6733 7644
rect 6789 7642 6813 7644
rect 6869 7642 6893 7644
rect 6949 7642 6973 7644
rect 7029 7642 7035 7644
rect 6789 7590 6791 7642
rect 6971 7590 6973 7642
rect 6727 7588 6733 7590
rect 6789 7588 6813 7590
rect 6869 7588 6893 7590
rect 6949 7588 6973 7590
rect 7029 7588 7035 7590
rect 6727 7579 7035 7588
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6656 6798 6684 7414
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7116 6662 7144 8502
rect 7300 6662 7328 8910
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7392 6848 7420 8842
rect 7484 7954 7512 9046
rect 7668 9030 7880 9058
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7472 6860 7524 6866
rect 7392 6820 7472 6848
rect 7472 6802 7524 6808
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 6727 6556 7035 6565
rect 6727 6554 6733 6556
rect 6789 6554 6813 6556
rect 6869 6554 6893 6556
rect 6949 6554 6973 6556
rect 7029 6554 7035 6556
rect 6789 6502 6791 6554
rect 6971 6502 6973 6554
rect 6727 6500 6733 6502
rect 6789 6500 6813 6502
rect 6869 6500 6893 6502
rect 6949 6500 6973 6502
rect 7029 6500 7035 6502
rect 6727 6491 7035 6500
rect 7300 6390 7328 6598
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6564 5681 6592 5782
rect 6550 5672 6606 5681
rect 6550 5607 6606 5616
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 5234 6684 5510
rect 6727 5468 7035 5477
rect 6727 5466 6733 5468
rect 6789 5466 6813 5468
rect 6869 5466 6893 5468
rect 6949 5466 6973 5468
rect 7029 5466 7035 5468
rect 6789 5414 6791 5466
rect 6971 5414 6973 5466
rect 6727 5412 6733 5414
rect 6789 5412 6813 5414
rect 6869 5412 6893 5414
rect 6949 5412 6973 5414
rect 7029 5412 7035 5414
rect 6727 5403 7035 5412
rect 7300 5234 7328 6326
rect 7484 6322 7512 6802
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7576 6458 7604 6666
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 5814 4720 5870 4729
rect 5814 4655 5870 4664
rect 5828 4282 5856 4655
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 6472 4214 6500 4762
rect 6727 4380 7035 4389
rect 6727 4378 6733 4380
rect 6789 4378 6813 4380
rect 6869 4378 6893 4380
rect 6949 4378 6973 4380
rect 7029 4378 7035 4380
rect 6789 4326 6791 4378
rect 6971 4326 6973 4378
rect 6727 4324 6733 4326
rect 6789 4324 6813 4326
rect 6869 4324 6893 4326
rect 6949 4324 6973 4326
rect 7029 4324 7035 4326
rect 6727 4315 7035 4324
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 5908 3936 5960 3942
rect 6380 3924 6408 4082
rect 6460 3936 6512 3942
rect 6380 3896 6460 3924
rect 5908 3878 5960 3884
rect 6460 3878 6512 3884
rect 5920 3738 5948 3878
rect 6067 3836 6375 3845
rect 6067 3834 6073 3836
rect 6129 3834 6153 3836
rect 6209 3834 6233 3836
rect 6289 3834 6313 3836
rect 6369 3834 6375 3836
rect 6129 3782 6131 3834
rect 6311 3782 6313 3834
rect 6067 3780 6073 3782
rect 6129 3780 6153 3782
rect 6209 3780 6233 3782
rect 6289 3780 6313 3782
rect 6369 3780 6375 3782
rect 6067 3771 6375 3780
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5262 2952 5318 2961
rect 5262 2887 5318 2896
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 3804 2746 3924 2774
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3528 2310 3556 2746
rect 3896 2446 3924 2746
rect 4020 2748 4328 2757
rect 4020 2746 4026 2748
rect 4082 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4328 2748
rect 4082 2694 4084 2746
rect 4264 2694 4266 2746
rect 4020 2692 4026 2694
rect 4082 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4328 2694
rect 4020 2683 4328 2692
rect 4448 2650 4476 2790
rect 5736 2774 5764 2994
rect 5920 2854 5948 3334
rect 6472 3194 6500 3878
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6564 3058 6592 3470
rect 6656 3194 6684 4218
rect 7300 4078 7328 5170
rect 7484 4622 7512 6258
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7576 5273 7604 5306
rect 7562 5264 7618 5273
rect 7562 5199 7618 5208
rect 7668 5166 7696 6734
rect 7760 6730 7788 9030
rect 8496 8634 8524 9930
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8588 9518 8616 9862
rect 8774 9820 9082 9829
rect 8774 9818 8780 9820
rect 8836 9818 8860 9820
rect 8916 9818 8940 9820
rect 8996 9818 9020 9820
rect 9076 9818 9082 9820
rect 8836 9766 8838 9818
rect 9018 9766 9020 9818
rect 8774 9764 8780 9766
rect 8836 9764 8860 9766
rect 8916 9764 8940 9766
rect 8996 9764 9020 9766
rect 9076 9764 9082 9766
rect 8774 9755 9082 9764
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8588 9110 8616 9454
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8774 8732 9082 8741
rect 8774 8730 8780 8732
rect 8836 8730 8860 8732
rect 8916 8730 8940 8732
rect 8996 8730 9020 8732
rect 9076 8730 9082 8732
rect 8836 8678 8838 8730
rect 9018 8678 9020 8730
rect 8774 8676 8780 8678
rect 8836 8676 8860 8678
rect 8916 8676 8940 8678
rect 8996 8676 9020 8678
rect 9076 8676 9082 8678
rect 8774 8667 9082 8676
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 9218 8256 9274 8265
rect 8114 8188 8422 8197
rect 9218 8191 9274 8200
rect 8114 8186 8120 8188
rect 8176 8186 8200 8188
rect 8256 8186 8280 8188
rect 8336 8186 8360 8188
rect 8416 8186 8422 8188
rect 8176 8134 8178 8186
rect 8358 8134 8360 8186
rect 8114 8132 8120 8134
rect 8176 8132 8200 8134
rect 8256 8132 8280 8134
rect 8336 8132 8360 8134
rect 8416 8132 8422 8134
rect 8114 8123 8422 8132
rect 9232 7886 9260 8191
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7852 7002 7880 7142
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7944 6934 7972 7142
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7748 6724 7800 6730
rect 7800 6684 7880 6712
rect 7748 6666 7800 6672
rect 7852 6322 7880 6684
rect 7944 6338 7972 6870
rect 8036 6866 8064 7414
rect 8114 7100 8422 7109
rect 8114 7098 8120 7100
rect 8176 7098 8200 7100
rect 8256 7098 8280 7100
rect 8336 7098 8360 7100
rect 8416 7098 8422 7100
rect 8176 7046 8178 7098
rect 8358 7046 8360 7098
rect 8114 7044 8120 7046
rect 8176 7044 8200 7046
rect 8256 7044 8280 7046
rect 8336 7044 8360 7046
rect 8416 7044 8422 7046
rect 8114 7035 8422 7044
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8036 6458 8064 6802
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7840 6316 7892 6322
rect 7944 6310 8064 6338
rect 7840 6258 7892 6264
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 6727 3292 7035 3301
rect 6727 3290 6733 3292
rect 6789 3290 6813 3292
rect 6869 3290 6893 3292
rect 6949 3290 6973 3292
rect 7029 3290 7035 3292
rect 6789 3238 6791 3290
rect 6971 3238 6973 3290
rect 6727 3236 6733 3238
rect 6789 3236 6813 3238
rect 6869 3236 6893 3238
rect 6949 3236 6973 3238
rect 7029 3236 7035 3238
rect 6727 3227 7035 3236
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5644 2746 5764 2774
rect 7760 2774 7788 6054
rect 7852 5846 7880 6258
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7944 5234 7972 6122
rect 8036 6118 8064 6310
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8114 6012 8422 6021
rect 8114 6010 8120 6012
rect 8176 6010 8200 6012
rect 8256 6010 8280 6012
rect 8336 6010 8360 6012
rect 8416 6010 8422 6012
rect 8176 5958 8178 6010
rect 8358 5958 8360 6010
rect 8114 5956 8120 5958
rect 8176 5956 8200 5958
rect 8256 5956 8280 5958
rect 8336 5956 8360 5958
rect 8416 5956 8422 5958
rect 8114 5947 8422 5956
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8496 5030 8524 7754
rect 8774 7644 9082 7653
rect 8774 7642 8780 7644
rect 8836 7642 8860 7644
rect 8916 7642 8940 7644
rect 8996 7642 9020 7644
rect 9076 7642 9082 7644
rect 8836 7590 8838 7642
rect 9018 7590 9020 7642
rect 8774 7588 8780 7590
rect 8836 7588 8860 7590
rect 8916 7588 8940 7590
rect 8996 7588 9020 7590
rect 9076 7588 9082 7590
rect 8774 7579 9082 7588
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8680 6798 8708 7414
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6322 8616 6598
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8114 4924 8422 4933
rect 8114 4922 8120 4924
rect 8176 4922 8200 4924
rect 8256 4922 8280 4924
rect 8336 4922 8360 4924
rect 8416 4922 8422 4924
rect 8176 4870 8178 4922
rect 8358 4870 8360 4922
rect 8114 4868 8120 4870
rect 8176 4868 8200 4870
rect 8256 4868 8280 4870
rect 8336 4868 8360 4870
rect 8416 4868 8422 4870
rect 8114 4859 8422 4868
rect 8496 4146 8524 4966
rect 8680 4554 8708 6734
rect 8774 6556 9082 6565
rect 8774 6554 8780 6556
rect 8836 6554 8860 6556
rect 8916 6554 8940 6556
rect 8996 6554 9020 6556
rect 9076 6554 9082 6556
rect 8836 6502 8838 6554
rect 9018 6502 9020 6554
rect 8774 6500 8780 6502
rect 8836 6500 8860 6502
rect 8916 6500 8940 6502
rect 8996 6500 9020 6502
rect 9076 6500 9082 6502
rect 8774 6491 9082 6500
rect 9312 5568 9364 5574
rect 9310 5536 9312 5545
rect 9364 5536 9366 5545
rect 8774 5468 9082 5477
rect 9310 5471 9366 5480
rect 8774 5466 8780 5468
rect 8836 5466 8860 5468
rect 8916 5466 8940 5468
rect 8996 5466 9020 5468
rect 9076 5466 9082 5468
rect 8836 5414 8838 5466
rect 9018 5414 9020 5466
rect 8774 5412 8780 5414
rect 8836 5412 8860 5414
rect 8916 5412 8940 5414
rect 8996 5412 9020 5414
rect 9076 5412 9082 5414
rect 8774 5403 9082 5412
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8114 3836 8422 3845
rect 8114 3834 8120 3836
rect 8176 3834 8200 3836
rect 8256 3834 8280 3836
rect 8336 3834 8360 3836
rect 8416 3834 8422 3836
rect 8176 3782 8178 3834
rect 8358 3782 8360 3834
rect 8114 3780 8120 3782
rect 8176 3780 8200 3782
rect 8256 3780 8280 3782
rect 8336 3780 8360 3782
rect 8416 3780 8422 3782
rect 8114 3771 8422 3780
rect 6067 2748 6375 2757
rect 6067 2746 6073 2748
rect 6129 2746 6153 2748
rect 6209 2746 6233 2748
rect 6289 2746 6313 2748
rect 6369 2746 6375 2748
rect 7760 2746 7880 2774
rect 5644 2650 5672 2746
rect 6129 2694 6131 2746
rect 6311 2694 6313 2746
rect 6067 2692 6073 2694
rect 6129 2692 6153 2694
rect 6209 2692 6233 2694
rect 6289 2692 6313 2694
rect 6369 2692 6375 2694
rect 6067 2683 6375 2692
rect 7852 2650 7880 2746
rect 8114 2748 8422 2757
rect 8114 2746 8120 2748
rect 8176 2746 8200 2748
rect 8256 2746 8280 2748
rect 8336 2746 8360 2748
rect 8416 2746 8422 2748
rect 8176 2694 8178 2746
rect 8358 2694 8360 2746
rect 8114 2692 8120 2694
rect 8176 2692 8200 2694
rect 8256 2692 8280 2694
rect 8336 2692 8360 2694
rect 8416 2692 8422 2694
rect 8114 2683 8422 2692
rect 8680 2650 8708 4490
rect 8774 4380 9082 4389
rect 8774 4378 8780 4380
rect 8836 4378 8860 4380
rect 8916 4378 8940 4380
rect 8996 4378 9020 4380
rect 9076 4378 9082 4380
rect 8836 4326 8838 4378
rect 9018 4326 9020 4378
rect 8774 4324 8780 4326
rect 8836 4324 8860 4326
rect 8916 4324 8940 4326
rect 8996 4324 9020 4326
rect 9076 4324 9082 4326
rect 8774 4315 9082 4324
rect 8774 3292 9082 3301
rect 8774 3290 8780 3292
rect 8836 3290 8860 3292
rect 8916 3290 8940 3292
rect 8996 3290 9020 3292
rect 9076 3290 9082 3292
rect 8836 3238 8838 3290
rect 9018 3238 9020 3290
rect 8774 3236 8780 3238
rect 8836 3236 8860 3238
rect 8916 3236 8940 3238
rect 8996 3236 9020 3238
rect 9076 3236 9082 3238
rect 8774 3227 9082 3236
rect 8852 2848 8904 2854
rect 8850 2816 8852 2825
rect 8904 2816 8906 2825
rect 8850 2751 8906 2760
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 2633 2204 2941 2213
rect 2633 2202 2639 2204
rect 2695 2202 2719 2204
rect 2775 2202 2799 2204
rect 2855 2202 2879 2204
rect 2935 2202 2941 2204
rect 2695 2150 2697 2202
rect 2877 2150 2879 2202
rect 2633 2148 2639 2150
rect 2695 2148 2719 2150
rect 2775 2148 2799 2150
rect 2855 2148 2879 2150
rect 2935 2148 2941 2150
rect 2633 2139 2941 2148
rect 4680 2204 4988 2213
rect 4680 2202 4686 2204
rect 4742 2202 4766 2204
rect 4822 2202 4846 2204
rect 4902 2202 4926 2204
rect 4982 2202 4988 2204
rect 4742 2150 4744 2202
rect 4924 2150 4926 2202
rect 4680 2148 4686 2150
rect 4742 2148 4766 2150
rect 4822 2148 4846 2150
rect 4902 2148 4926 2150
rect 4982 2148 4988 2150
rect 4680 2139 4988 2148
rect 2516 1958 2636 1986
rect 2608 800 2636 1958
rect 5276 1306 5304 2382
rect 6727 2204 7035 2213
rect 6727 2202 6733 2204
rect 6789 2202 6813 2204
rect 6869 2202 6893 2204
rect 6949 2202 6973 2204
rect 7029 2202 7035 2204
rect 6789 2150 6791 2202
rect 6971 2150 6973 2202
rect 6727 2148 6733 2150
rect 6789 2148 6813 2150
rect 6869 2148 6893 2150
rect 6949 2148 6973 2150
rect 7029 2148 7035 2150
rect 6727 2139 7035 2148
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 7760 800 7788 2382
rect 8774 2204 9082 2213
rect 8774 2202 8780 2204
rect 8836 2202 8860 2204
rect 8916 2202 8940 2204
rect 8996 2202 9020 2204
rect 9076 2202 9082 2204
rect 8836 2150 8838 2202
rect 9018 2150 9020 2202
rect 8774 2148 8780 2150
rect 8836 2148 8860 2150
rect 8916 2148 8940 2150
rect 8996 2148 9020 2150
rect 9076 2148 9082 2150
rect 8774 2139 9082 2148
rect 10336 800 10364 2382
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 7746 0 7802 800
rect 10322 0 10378 800
<< via2 >>
rect 938 10920 994 10976
rect 1979 10362 2035 10364
rect 2059 10362 2115 10364
rect 2139 10362 2195 10364
rect 2219 10362 2275 10364
rect 1979 10310 2025 10362
rect 2025 10310 2035 10362
rect 2059 10310 2089 10362
rect 2089 10310 2101 10362
rect 2101 10310 2115 10362
rect 2139 10310 2153 10362
rect 2153 10310 2165 10362
rect 2165 10310 2195 10362
rect 2219 10310 2229 10362
rect 2229 10310 2275 10362
rect 1979 10308 2035 10310
rect 2059 10308 2115 10310
rect 2139 10308 2195 10310
rect 2219 10308 2275 10310
rect 1398 8200 1454 8256
rect 2639 9818 2695 9820
rect 2719 9818 2775 9820
rect 2799 9818 2855 9820
rect 2879 9818 2935 9820
rect 2639 9766 2685 9818
rect 2685 9766 2695 9818
rect 2719 9766 2749 9818
rect 2749 9766 2761 9818
rect 2761 9766 2775 9818
rect 2799 9766 2813 9818
rect 2813 9766 2825 9818
rect 2825 9766 2855 9818
rect 2879 9766 2889 9818
rect 2889 9766 2935 9818
rect 2639 9764 2695 9766
rect 2719 9764 2775 9766
rect 2799 9764 2855 9766
rect 2879 9764 2935 9766
rect 4026 10362 4082 10364
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4026 10310 4072 10362
rect 4072 10310 4082 10362
rect 4106 10310 4136 10362
rect 4136 10310 4148 10362
rect 4148 10310 4162 10362
rect 4186 10310 4200 10362
rect 4200 10310 4212 10362
rect 4212 10310 4242 10362
rect 4266 10310 4276 10362
rect 4276 10310 4322 10362
rect 4026 10308 4082 10310
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 6073 10362 6129 10364
rect 6153 10362 6209 10364
rect 6233 10362 6289 10364
rect 6313 10362 6369 10364
rect 6073 10310 6119 10362
rect 6119 10310 6129 10362
rect 6153 10310 6183 10362
rect 6183 10310 6195 10362
rect 6195 10310 6209 10362
rect 6233 10310 6247 10362
rect 6247 10310 6259 10362
rect 6259 10310 6289 10362
rect 6313 10310 6323 10362
rect 6323 10310 6369 10362
rect 6073 10308 6129 10310
rect 6153 10308 6209 10310
rect 6233 10308 6289 10310
rect 6313 10308 6369 10310
rect 8120 10362 8176 10364
rect 8200 10362 8256 10364
rect 8280 10362 8336 10364
rect 8360 10362 8416 10364
rect 8120 10310 8166 10362
rect 8166 10310 8176 10362
rect 8200 10310 8230 10362
rect 8230 10310 8242 10362
rect 8242 10310 8256 10362
rect 8280 10310 8294 10362
rect 8294 10310 8306 10362
rect 8306 10310 8336 10362
rect 8360 10310 8370 10362
rect 8370 10310 8416 10362
rect 8120 10308 8176 10310
rect 8200 10308 8256 10310
rect 8280 10308 8336 10310
rect 8360 10308 8416 10310
rect 9218 10920 9274 10976
rect 4686 9818 4742 9820
rect 4766 9818 4822 9820
rect 4846 9818 4902 9820
rect 4926 9818 4982 9820
rect 4686 9766 4732 9818
rect 4732 9766 4742 9818
rect 4766 9766 4796 9818
rect 4796 9766 4808 9818
rect 4808 9766 4822 9818
rect 4846 9766 4860 9818
rect 4860 9766 4872 9818
rect 4872 9766 4902 9818
rect 4926 9766 4936 9818
rect 4936 9766 4982 9818
rect 4686 9764 4742 9766
rect 4766 9764 4822 9766
rect 4846 9764 4902 9766
rect 4926 9764 4982 9766
rect 1979 9274 2035 9276
rect 2059 9274 2115 9276
rect 2139 9274 2195 9276
rect 2219 9274 2275 9276
rect 1979 9222 2025 9274
rect 2025 9222 2035 9274
rect 2059 9222 2089 9274
rect 2089 9222 2101 9274
rect 2101 9222 2115 9274
rect 2139 9222 2153 9274
rect 2153 9222 2165 9274
rect 2165 9222 2195 9274
rect 2219 9222 2229 9274
rect 2229 9222 2275 9274
rect 1979 9220 2035 9222
rect 2059 9220 2115 9222
rect 2139 9220 2195 9222
rect 2219 9220 2275 9222
rect 2639 8730 2695 8732
rect 2719 8730 2775 8732
rect 2799 8730 2855 8732
rect 2879 8730 2935 8732
rect 2639 8678 2685 8730
rect 2685 8678 2695 8730
rect 2719 8678 2749 8730
rect 2749 8678 2761 8730
rect 2761 8678 2775 8730
rect 2799 8678 2813 8730
rect 2813 8678 2825 8730
rect 2825 8678 2855 8730
rect 2879 8678 2889 8730
rect 2889 8678 2935 8730
rect 2639 8676 2695 8678
rect 2719 8676 2775 8678
rect 2799 8676 2855 8678
rect 2879 8676 2935 8678
rect 1979 8186 2035 8188
rect 2059 8186 2115 8188
rect 2139 8186 2195 8188
rect 2219 8186 2275 8188
rect 1979 8134 2025 8186
rect 2025 8134 2035 8186
rect 2059 8134 2089 8186
rect 2089 8134 2101 8186
rect 2101 8134 2115 8186
rect 2139 8134 2153 8186
rect 2153 8134 2165 8186
rect 2165 8134 2195 8186
rect 2219 8134 2229 8186
rect 2229 8134 2275 8186
rect 1979 8132 2035 8134
rect 2059 8132 2115 8134
rect 2139 8132 2195 8134
rect 2219 8132 2275 8134
rect 2639 7642 2695 7644
rect 2719 7642 2775 7644
rect 2799 7642 2855 7644
rect 2879 7642 2935 7644
rect 2639 7590 2685 7642
rect 2685 7590 2695 7642
rect 2719 7590 2749 7642
rect 2749 7590 2761 7642
rect 2761 7590 2775 7642
rect 2799 7590 2813 7642
rect 2813 7590 2825 7642
rect 2825 7590 2855 7642
rect 2879 7590 2889 7642
rect 2889 7590 2935 7642
rect 2639 7588 2695 7590
rect 2719 7588 2775 7590
rect 2799 7588 2855 7590
rect 2879 7588 2935 7590
rect 1979 7098 2035 7100
rect 2059 7098 2115 7100
rect 2139 7098 2195 7100
rect 2219 7098 2275 7100
rect 1979 7046 2025 7098
rect 2025 7046 2035 7098
rect 2059 7046 2089 7098
rect 2089 7046 2101 7098
rect 2101 7046 2115 7098
rect 2139 7046 2153 7098
rect 2153 7046 2165 7098
rect 2165 7046 2195 7098
rect 2219 7046 2229 7098
rect 2229 7046 2275 7098
rect 1979 7044 2035 7046
rect 2059 7044 2115 7046
rect 2139 7044 2195 7046
rect 2219 7044 2275 7046
rect 2639 6554 2695 6556
rect 2719 6554 2775 6556
rect 2799 6554 2855 6556
rect 2879 6554 2935 6556
rect 2639 6502 2685 6554
rect 2685 6502 2695 6554
rect 2719 6502 2749 6554
rect 2749 6502 2761 6554
rect 2761 6502 2775 6554
rect 2799 6502 2813 6554
rect 2813 6502 2825 6554
rect 2825 6502 2855 6554
rect 2879 6502 2889 6554
rect 2889 6502 2935 6554
rect 2639 6500 2695 6502
rect 2719 6500 2775 6502
rect 2799 6500 2855 6502
rect 2879 6500 2935 6502
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 1582 5480 1638 5516
rect 1979 6010 2035 6012
rect 2059 6010 2115 6012
rect 2139 6010 2195 6012
rect 2219 6010 2275 6012
rect 1979 5958 2025 6010
rect 2025 5958 2035 6010
rect 2059 5958 2089 6010
rect 2089 5958 2101 6010
rect 2101 5958 2115 6010
rect 2139 5958 2153 6010
rect 2153 5958 2165 6010
rect 2165 5958 2195 6010
rect 2219 5958 2229 6010
rect 2229 5958 2275 6010
rect 1979 5956 2035 5958
rect 2059 5956 2115 5958
rect 2139 5956 2195 5958
rect 2219 5956 2275 5958
rect 2639 5466 2695 5468
rect 2719 5466 2775 5468
rect 2799 5466 2855 5468
rect 2879 5466 2935 5468
rect 2639 5414 2685 5466
rect 2685 5414 2695 5466
rect 2719 5414 2749 5466
rect 2749 5414 2761 5466
rect 2761 5414 2775 5466
rect 2799 5414 2813 5466
rect 2813 5414 2825 5466
rect 2825 5414 2855 5466
rect 2879 5414 2889 5466
rect 2889 5414 2935 5466
rect 2639 5412 2695 5414
rect 2719 5412 2775 5414
rect 2799 5412 2855 5414
rect 2879 5412 2935 5414
rect 4026 9274 4082 9276
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4026 9222 4072 9274
rect 4072 9222 4082 9274
rect 4106 9222 4136 9274
rect 4136 9222 4148 9274
rect 4148 9222 4162 9274
rect 4186 9222 4200 9274
rect 4200 9222 4212 9274
rect 4212 9222 4242 9274
rect 4266 9222 4276 9274
rect 4276 9222 4322 9274
rect 4026 9220 4082 9222
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 4686 8730 4742 8732
rect 4766 8730 4822 8732
rect 4846 8730 4902 8732
rect 4926 8730 4982 8732
rect 4686 8678 4732 8730
rect 4732 8678 4742 8730
rect 4766 8678 4796 8730
rect 4796 8678 4808 8730
rect 4808 8678 4822 8730
rect 4846 8678 4860 8730
rect 4860 8678 4872 8730
rect 4872 8678 4902 8730
rect 4926 8678 4936 8730
rect 4936 8678 4982 8730
rect 4686 8676 4742 8678
rect 4766 8676 4822 8678
rect 4846 8676 4902 8678
rect 4926 8676 4982 8678
rect 4026 8186 4082 8188
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4026 8134 4072 8186
rect 4072 8134 4082 8186
rect 4106 8134 4136 8186
rect 4136 8134 4148 8186
rect 4148 8134 4162 8186
rect 4186 8134 4200 8186
rect 4200 8134 4212 8186
rect 4212 8134 4242 8186
rect 4266 8134 4276 8186
rect 4276 8134 4322 8186
rect 4026 8132 4082 8134
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 1979 4922 2035 4924
rect 2059 4922 2115 4924
rect 2139 4922 2195 4924
rect 2219 4922 2275 4924
rect 1979 4870 2025 4922
rect 2025 4870 2035 4922
rect 2059 4870 2089 4922
rect 2089 4870 2101 4922
rect 2101 4870 2115 4922
rect 2139 4870 2153 4922
rect 2153 4870 2165 4922
rect 2165 4870 2195 4922
rect 2219 4870 2229 4922
rect 2229 4870 2275 4922
rect 1979 4868 2035 4870
rect 2059 4868 2115 4870
rect 2139 4868 2195 4870
rect 2219 4868 2275 4870
rect 1979 3834 2035 3836
rect 2059 3834 2115 3836
rect 2139 3834 2195 3836
rect 2219 3834 2275 3836
rect 1979 3782 2025 3834
rect 2025 3782 2035 3834
rect 2059 3782 2089 3834
rect 2089 3782 2101 3834
rect 2101 3782 2115 3834
rect 2139 3782 2153 3834
rect 2153 3782 2165 3834
rect 2165 3782 2195 3834
rect 2219 3782 2229 3834
rect 2229 3782 2275 3834
rect 1979 3780 2035 3782
rect 2059 3780 2115 3782
rect 2139 3780 2195 3782
rect 2219 3780 2275 3782
rect 2639 4378 2695 4380
rect 2719 4378 2775 4380
rect 2799 4378 2855 4380
rect 2879 4378 2935 4380
rect 2639 4326 2685 4378
rect 2685 4326 2695 4378
rect 2719 4326 2749 4378
rect 2749 4326 2761 4378
rect 2761 4326 2775 4378
rect 2799 4326 2813 4378
rect 2813 4326 2825 4378
rect 2825 4326 2855 4378
rect 2879 4326 2889 4378
rect 2889 4326 2935 4378
rect 2639 4324 2695 4326
rect 2719 4324 2775 4326
rect 2799 4324 2855 4326
rect 2879 4324 2935 4326
rect 938 2760 994 2816
rect 2639 3290 2695 3292
rect 2719 3290 2775 3292
rect 2799 3290 2855 3292
rect 2879 3290 2935 3292
rect 2639 3238 2685 3290
rect 2685 3238 2695 3290
rect 2719 3238 2749 3290
rect 2749 3238 2761 3290
rect 2761 3238 2775 3290
rect 2799 3238 2813 3290
rect 2813 3238 2825 3290
rect 2825 3238 2855 3290
rect 2879 3238 2889 3290
rect 2889 3238 2935 3290
rect 2639 3236 2695 3238
rect 2719 3236 2775 3238
rect 2799 3236 2855 3238
rect 2879 3236 2935 3238
rect 2502 2896 2558 2952
rect 1979 2746 2035 2748
rect 2059 2746 2115 2748
rect 2139 2746 2195 2748
rect 2219 2746 2275 2748
rect 1979 2694 2025 2746
rect 2025 2694 2035 2746
rect 2059 2694 2089 2746
rect 2089 2694 2101 2746
rect 2101 2694 2115 2746
rect 2139 2694 2153 2746
rect 2153 2694 2165 2746
rect 2165 2694 2195 2746
rect 2219 2694 2229 2746
rect 2229 2694 2275 2746
rect 1979 2692 2035 2694
rect 2059 2692 2115 2694
rect 2139 2692 2195 2694
rect 2219 2692 2275 2694
rect 4686 7642 4742 7644
rect 4766 7642 4822 7644
rect 4846 7642 4902 7644
rect 4926 7642 4982 7644
rect 4686 7590 4732 7642
rect 4732 7590 4742 7642
rect 4766 7590 4796 7642
rect 4796 7590 4808 7642
rect 4808 7590 4822 7642
rect 4846 7590 4860 7642
rect 4860 7590 4872 7642
rect 4872 7590 4902 7642
rect 4926 7590 4936 7642
rect 4936 7590 4982 7642
rect 4686 7588 4742 7590
rect 4766 7588 4822 7590
rect 4846 7588 4902 7590
rect 4926 7588 4982 7590
rect 4026 7098 4082 7100
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4026 7046 4072 7098
rect 4072 7046 4082 7098
rect 4106 7046 4136 7098
rect 4136 7046 4148 7098
rect 4148 7046 4162 7098
rect 4186 7046 4200 7098
rect 4200 7046 4212 7098
rect 4212 7046 4242 7098
rect 4266 7046 4276 7098
rect 4276 7046 4322 7098
rect 4026 7044 4082 7046
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 4026 6010 4082 6012
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4026 5958 4072 6010
rect 4072 5958 4082 6010
rect 4106 5958 4136 6010
rect 4136 5958 4148 6010
rect 4148 5958 4162 6010
rect 4186 5958 4200 6010
rect 4200 5958 4212 6010
rect 4212 5958 4242 6010
rect 4266 5958 4276 6010
rect 4276 5958 4322 6010
rect 4026 5956 4082 5958
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4158 5752 4214 5808
rect 4686 6554 4742 6556
rect 4766 6554 4822 6556
rect 4846 6554 4902 6556
rect 4926 6554 4982 6556
rect 4686 6502 4732 6554
rect 4732 6502 4742 6554
rect 4766 6502 4796 6554
rect 4796 6502 4808 6554
rect 4808 6502 4822 6554
rect 4846 6502 4860 6554
rect 4860 6502 4872 6554
rect 4872 6502 4902 6554
rect 4926 6502 4936 6554
rect 4936 6502 4982 6554
rect 4686 6500 4742 6502
rect 4766 6500 4822 6502
rect 4846 6500 4902 6502
rect 4926 6500 4982 6502
rect 4342 5616 4398 5672
rect 4026 4922 4082 4924
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4026 4870 4072 4922
rect 4072 4870 4082 4922
rect 4106 4870 4136 4922
rect 4136 4870 4148 4922
rect 4148 4870 4162 4922
rect 4186 4870 4200 4922
rect 4200 4870 4212 4922
rect 4212 4870 4242 4922
rect 4266 4870 4276 4922
rect 4276 4870 4322 4922
rect 4026 4868 4082 4870
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4026 3834 4082 3836
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4026 3782 4072 3834
rect 4072 3782 4082 3834
rect 4106 3782 4136 3834
rect 4136 3782 4148 3834
rect 4148 3782 4162 3834
rect 4186 3782 4200 3834
rect 4200 3782 4212 3834
rect 4212 3782 4242 3834
rect 4266 3782 4276 3834
rect 4276 3782 4322 3834
rect 4026 3780 4082 3782
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4686 5466 4742 5468
rect 4766 5466 4822 5468
rect 4846 5466 4902 5468
rect 4926 5466 4982 5468
rect 4686 5414 4732 5466
rect 4732 5414 4742 5466
rect 4766 5414 4796 5466
rect 4796 5414 4808 5466
rect 4808 5414 4822 5466
rect 4846 5414 4860 5466
rect 4860 5414 4872 5466
rect 4872 5414 4902 5466
rect 4926 5414 4936 5466
rect 4936 5414 4982 5466
rect 4686 5412 4742 5414
rect 4766 5412 4822 5414
rect 4846 5412 4902 5414
rect 4926 5412 4982 5414
rect 4894 5228 4950 5264
rect 4894 5208 4896 5228
rect 4896 5208 4948 5228
rect 4948 5208 4950 5228
rect 5170 4664 5226 4720
rect 4686 4378 4742 4380
rect 4766 4378 4822 4380
rect 4846 4378 4902 4380
rect 4926 4378 4982 4380
rect 4686 4326 4732 4378
rect 4732 4326 4742 4378
rect 4766 4326 4796 4378
rect 4796 4326 4808 4378
rect 4808 4326 4822 4378
rect 4846 4326 4860 4378
rect 4860 4326 4872 4378
rect 4872 4326 4902 4378
rect 4926 4326 4936 4378
rect 4936 4326 4982 4378
rect 4686 4324 4742 4326
rect 4766 4324 4822 4326
rect 4846 4324 4902 4326
rect 4926 4324 4982 4326
rect 4686 3290 4742 3292
rect 4766 3290 4822 3292
rect 4846 3290 4902 3292
rect 4926 3290 4982 3292
rect 4686 3238 4732 3290
rect 4732 3238 4742 3290
rect 4766 3238 4796 3290
rect 4796 3238 4808 3290
rect 4808 3238 4822 3290
rect 4846 3238 4860 3290
rect 4860 3238 4872 3290
rect 4872 3238 4902 3290
rect 4926 3238 4936 3290
rect 4936 3238 4982 3290
rect 4686 3236 4742 3238
rect 4766 3236 4822 3238
rect 4846 3236 4902 3238
rect 4926 3236 4982 3238
rect 5446 5752 5502 5808
rect 6073 9274 6129 9276
rect 6153 9274 6209 9276
rect 6233 9274 6289 9276
rect 6313 9274 6369 9276
rect 6073 9222 6119 9274
rect 6119 9222 6129 9274
rect 6153 9222 6183 9274
rect 6183 9222 6195 9274
rect 6195 9222 6209 9274
rect 6233 9222 6247 9274
rect 6247 9222 6259 9274
rect 6259 9222 6289 9274
rect 6313 9222 6323 9274
rect 6323 9222 6369 9274
rect 6073 9220 6129 9222
rect 6153 9220 6209 9222
rect 6233 9220 6289 9222
rect 6313 9220 6369 9222
rect 6073 8186 6129 8188
rect 6153 8186 6209 8188
rect 6233 8186 6289 8188
rect 6313 8186 6369 8188
rect 6073 8134 6119 8186
rect 6119 8134 6129 8186
rect 6153 8134 6183 8186
rect 6183 8134 6195 8186
rect 6195 8134 6209 8186
rect 6233 8134 6247 8186
rect 6247 8134 6259 8186
rect 6259 8134 6289 8186
rect 6313 8134 6323 8186
rect 6323 8134 6369 8186
rect 6073 8132 6129 8134
rect 6153 8132 6209 8134
rect 6233 8132 6289 8134
rect 6313 8132 6369 8134
rect 6073 7098 6129 7100
rect 6153 7098 6209 7100
rect 6233 7098 6289 7100
rect 6313 7098 6369 7100
rect 6073 7046 6119 7098
rect 6119 7046 6129 7098
rect 6153 7046 6183 7098
rect 6183 7046 6195 7098
rect 6195 7046 6209 7098
rect 6233 7046 6247 7098
rect 6247 7046 6259 7098
rect 6259 7046 6289 7098
rect 6313 7046 6323 7098
rect 6323 7046 6369 7098
rect 6073 7044 6129 7046
rect 6153 7044 6209 7046
rect 6233 7044 6289 7046
rect 6313 7044 6369 7046
rect 6073 6010 6129 6012
rect 6153 6010 6209 6012
rect 6233 6010 6289 6012
rect 6313 6010 6369 6012
rect 6073 5958 6119 6010
rect 6119 5958 6129 6010
rect 6153 5958 6183 6010
rect 6183 5958 6195 6010
rect 6195 5958 6209 6010
rect 6233 5958 6247 6010
rect 6247 5958 6259 6010
rect 6259 5958 6289 6010
rect 6313 5958 6323 6010
rect 6323 5958 6369 6010
rect 6073 5956 6129 5958
rect 6153 5956 6209 5958
rect 6233 5956 6289 5958
rect 6313 5956 6369 5958
rect 6073 4922 6129 4924
rect 6153 4922 6209 4924
rect 6233 4922 6289 4924
rect 6313 4922 6369 4924
rect 6073 4870 6119 4922
rect 6119 4870 6129 4922
rect 6153 4870 6183 4922
rect 6183 4870 6195 4922
rect 6195 4870 6209 4922
rect 6233 4870 6247 4922
rect 6247 4870 6259 4922
rect 6259 4870 6289 4922
rect 6313 4870 6323 4922
rect 6323 4870 6369 4922
rect 6073 4868 6129 4870
rect 6153 4868 6209 4870
rect 6233 4868 6289 4870
rect 6313 4868 6369 4870
rect 6733 9818 6789 9820
rect 6813 9818 6869 9820
rect 6893 9818 6949 9820
rect 6973 9818 7029 9820
rect 6733 9766 6779 9818
rect 6779 9766 6789 9818
rect 6813 9766 6843 9818
rect 6843 9766 6855 9818
rect 6855 9766 6869 9818
rect 6893 9766 6907 9818
rect 6907 9766 6919 9818
rect 6919 9766 6949 9818
rect 6973 9766 6983 9818
rect 6983 9766 7029 9818
rect 6733 9764 6789 9766
rect 6813 9764 6869 9766
rect 6893 9764 6949 9766
rect 6973 9764 7029 9766
rect 8120 9274 8176 9276
rect 8200 9274 8256 9276
rect 8280 9274 8336 9276
rect 8360 9274 8416 9276
rect 8120 9222 8166 9274
rect 8166 9222 8176 9274
rect 8200 9222 8230 9274
rect 8230 9222 8242 9274
rect 8242 9222 8256 9274
rect 8280 9222 8294 9274
rect 8294 9222 8306 9274
rect 8306 9222 8336 9274
rect 8360 9222 8370 9274
rect 8370 9222 8416 9274
rect 8120 9220 8176 9222
rect 8200 9220 8256 9222
rect 8280 9220 8336 9222
rect 8360 9220 8416 9222
rect 6733 8730 6789 8732
rect 6813 8730 6869 8732
rect 6893 8730 6949 8732
rect 6973 8730 7029 8732
rect 6733 8678 6779 8730
rect 6779 8678 6789 8730
rect 6813 8678 6843 8730
rect 6843 8678 6855 8730
rect 6855 8678 6869 8730
rect 6893 8678 6907 8730
rect 6907 8678 6919 8730
rect 6919 8678 6949 8730
rect 6973 8678 6983 8730
rect 6983 8678 7029 8730
rect 6733 8676 6789 8678
rect 6813 8676 6869 8678
rect 6893 8676 6949 8678
rect 6973 8676 7029 8678
rect 6733 7642 6789 7644
rect 6813 7642 6869 7644
rect 6893 7642 6949 7644
rect 6973 7642 7029 7644
rect 6733 7590 6779 7642
rect 6779 7590 6789 7642
rect 6813 7590 6843 7642
rect 6843 7590 6855 7642
rect 6855 7590 6869 7642
rect 6893 7590 6907 7642
rect 6907 7590 6919 7642
rect 6919 7590 6949 7642
rect 6973 7590 6983 7642
rect 6983 7590 7029 7642
rect 6733 7588 6789 7590
rect 6813 7588 6869 7590
rect 6893 7588 6949 7590
rect 6973 7588 7029 7590
rect 6733 6554 6789 6556
rect 6813 6554 6869 6556
rect 6893 6554 6949 6556
rect 6973 6554 7029 6556
rect 6733 6502 6779 6554
rect 6779 6502 6789 6554
rect 6813 6502 6843 6554
rect 6843 6502 6855 6554
rect 6855 6502 6869 6554
rect 6893 6502 6907 6554
rect 6907 6502 6919 6554
rect 6919 6502 6949 6554
rect 6973 6502 6983 6554
rect 6983 6502 7029 6554
rect 6733 6500 6789 6502
rect 6813 6500 6869 6502
rect 6893 6500 6949 6502
rect 6973 6500 7029 6502
rect 6550 5616 6606 5672
rect 6733 5466 6789 5468
rect 6813 5466 6869 5468
rect 6893 5466 6949 5468
rect 6973 5466 7029 5468
rect 6733 5414 6779 5466
rect 6779 5414 6789 5466
rect 6813 5414 6843 5466
rect 6843 5414 6855 5466
rect 6855 5414 6869 5466
rect 6893 5414 6907 5466
rect 6907 5414 6919 5466
rect 6919 5414 6949 5466
rect 6973 5414 6983 5466
rect 6983 5414 7029 5466
rect 6733 5412 6789 5414
rect 6813 5412 6869 5414
rect 6893 5412 6949 5414
rect 6973 5412 7029 5414
rect 5814 4664 5870 4720
rect 6733 4378 6789 4380
rect 6813 4378 6869 4380
rect 6893 4378 6949 4380
rect 6973 4378 7029 4380
rect 6733 4326 6779 4378
rect 6779 4326 6789 4378
rect 6813 4326 6843 4378
rect 6843 4326 6855 4378
rect 6855 4326 6869 4378
rect 6893 4326 6907 4378
rect 6907 4326 6919 4378
rect 6919 4326 6949 4378
rect 6973 4326 6983 4378
rect 6983 4326 7029 4378
rect 6733 4324 6789 4326
rect 6813 4324 6869 4326
rect 6893 4324 6949 4326
rect 6973 4324 7029 4326
rect 6073 3834 6129 3836
rect 6153 3834 6209 3836
rect 6233 3834 6289 3836
rect 6313 3834 6369 3836
rect 6073 3782 6119 3834
rect 6119 3782 6129 3834
rect 6153 3782 6183 3834
rect 6183 3782 6195 3834
rect 6195 3782 6209 3834
rect 6233 3782 6247 3834
rect 6247 3782 6259 3834
rect 6259 3782 6289 3834
rect 6313 3782 6323 3834
rect 6323 3782 6369 3834
rect 6073 3780 6129 3782
rect 6153 3780 6209 3782
rect 6233 3780 6289 3782
rect 6313 3780 6369 3782
rect 5262 2896 5318 2952
rect 4026 2746 4082 2748
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4026 2694 4072 2746
rect 4072 2694 4082 2746
rect 4106 2694 4136 2746
rect 4136 2694 4148 2746
rect 4148 2694 4162 2746
rect 4186 2694 4200 2746
rect 4200 2694 4212 2746
rect 4212 2694 4242 2746
rect 4266 2694 4276 2746
rect 4276 2694 4322 2746
rect 4026 2692 4082 2694
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 7562 5208 7618 5264
rect 8780 9818 8836 9820
rect 8860 9818 8916 9820
rect 8940 9818 8996 9820
rect 9020 9818 9076 9820
rect 8780 9766 8826 9818
rect 8826 9766 8836 9818
rect 8860 9766 8890 9818
rect 8890 9766 8902 9818
rect 8902 9766 8916 9818
rect 8940 9766 8954 9818
rect 8954 9766 8966 9818
rect 8966 9766 8996 9818
rect 9020 9766 9030 9818
rect 9030 9766 9076 9818
rect 8780 9764 8836 9766
rect 8860 9764 8916 9766
rect 8940 9764 8996 9766
rect 9020 9764 9076 9766
rect 8780 8730 8836 8732
rect 8860 8730 8916 8732
rect 8940 8730 8996 8732
rect 9020 8730 9076 8732
rect 8780 8678 8826 8730
rect 8826 8678 8836 8730
rect 8860 8678 8890 8730
rect 8890 8678 8902 8730
rect 8902 8678 8916 8730
rect 8940 8678 8954 8730
rect 8954 8678 8966 8730
rect 8966 8678 8996 8730
rect 9020 8678 9030 8730
rect 9030 8678 9076 8730
rect 8780 8676 8836 8678
rect 8860 8676 8916 8678
rect 8940 8676 8996 8678
rect 9020 8676 9076 8678
rect 9218 8200 9274 8256
rect 8120 8186 8176 8188
rect 8200 8186 8256 8188
rect 8280 8186 8336 8188
rect 8360 8186 8416 8188
rect 8120 8134 8166 8186
rect 8166 8134 8176 8186
rect 8200 8134 8230 8186
rect 8230 8134 8242 8186
rect 8242 8134 8256 8186
rect 8280 8134 8294 8186
rect 8294 8134 8306 8186
rect 8306 8134 8336 8186
rect 8360 8134 8370 8186
rect 8370 8134 8416 8186
rect 8120 8132 8176 8134
rect 8200 8132 8256 8134
rect 8280 8132 8336 8134
rect 8360 8132 8416 8134
rect 8120 7098 8176 7100
rect 8200 7098 8256 7100
rect 8280 7098 8336 7100
rect 8360 7098 8416 7100
rect 8120 7046 8166 7098
rect 8166 7046 8176 7098
rect 8200 7046 8230 7098
rect 8230 7046 8242 7098
rect 8242 7046 8256 7098
rect 8280 7046 8294 7098
rect 8294 7046 8306 7098
rect 8306 7046 8336 7098
rect 8360 7046 8370 7098
rect 8370 7046 8416 7098
rect 8120 7044 8176 7046
rect 8200 7044 8256 7046
rect 8280 7044 8336 7046
rect 8360 7044 8416 7046
rect 6733 3290 6789 3292
rect 6813 3290 6869 3292
rect 6893 3290 6949 3292
rect 6973 3290 7029 3292
rect 6733 3238 6779 3290
rect 6779 3238 6789 3290
rect 6813 3238 6843 3290
rect 6843 3238 6855 3290
rect 6855 3238 6869 3290
rect 6893 3238 6907 3290
rect 6907 3238 6919 3290
rect 6919 3238 6949 3290
rect 6973 3238 6983 3290
rect 6983 3238 7029 3290
rect 6733 3236 6789 3238
rect 6813 3236 6869 3238
rect 6893 3236 6949 3238
rect 6973 3236 7029 3238
rect 8120 6010 8176 6012
rect 8200 6010 8256 6012
rect 8280 6010 8336 6012
rect 8360 6010 8416 6012
rect 8120 5958 8166 6010
rect 8166 5958 8176 6010
rect 8200 5958 8230 6010
rect 8230 5958 8242 6010
rect 8242 5958 8256 6010
rect 8280 5958 8294 6010
rect 8294 5958 8306 6010
rect 8306 5958 8336 6010
rect 8360 5958 8370 6010
rect 8370 5958 8416 6010
rect 8120 5956 8176 5958
rect 8200 5956 8256 5958
rect 8280 5956 8336 5958
rect 8360 5956 8416 5958
rect 8780 7642 8836 7644
rect 8860 7642 8916 7644
rect 8940 7642 8996 7644
rect 9020 7642 9076 7644
rect 8780 7590 8826 7642
rect 8826 7590 8836 7642
rect 8860 7590 8890 7642
rect 8890 7590 8902 7642
rect 8902 7590 8916 7642
rect 8940 7590 8954 7642
rect 8954 7590 8966 7642
rect 8966 7590 8996 7642
rect 9020 7590 9030 7642
rect 9030 7590 9076 7642
rect 8780 7588 8836 7590
rect 8860 7588 8916 7590
rect 8940 7588 8996 7590
rect 9020 7588 9076 7590
rect 8120 4922 8176 4924
rect 8200 4922 8256 4924
rect 8280 4922 8336 4924
rect 8360 4922 8416 4924
rect 8120 4870 8166 4922
rect 8166 4870 8176 4922
rect 8200 4870 8230 4922
rect 8230 4870 8242 4922
rect 8242 4870 8256 4922
rect 8280 4870 8294 4922
rect 8294 4870 8306 4922
rect 8306 4870 8336 4922
rect 8360 4870 8370 4922
rect 8370 4870 8416 4922
rect 8120 4868 8176 4870
rect 8200 4868 8256 4870
rect 8280 4868 8336 4870
rect 8360 4868 8416 4870
rect 8780 6554 8836 6556
rect 8860 6554 8916 6556
rect 8940 6554 8996 6556
rect 9020 6554 9076 6556
rect 8780 6502 8826 6554
rect 8826 6502 8836 6554
rect 8860 6502 8890 6554
rect 8890 6502 8902 6554
rect 8902 6502 8916 6554
rect 8940 6502 8954 6554
rect 8954 6502 8966 6554
rect 8966 6502 8996 6554
rect 9020 6502 9030 6554
rect 9030 6502 9076 6554
rect 8780 6500 8836 6502
rect 8860 6500 8916 6502
rect 8940 6500 8996 6502
rect 9020 6500 9076 6502
rect 9310 5516 9312 5536
rect 9312 5516 9364 5536
rect 9364 5516 9366 5536
rect 9310 5480 9366 5516
rect 8780 5466 8836 5468
rect 8860 5466 8916 5468
rect 8940 5466 8996 5468
rect 9020 5466 9076 5468
rect 8780 5414 8826 5466
rect 8826 5414 8836 5466
rect 8860 5414 8890 5466
rect 8890 5414 8902 5466
rect 8902 5414 8916 5466
rect 8940 5414 8954 5466
rect 8954 5414 8966 5466
rect 8966 5414 8996 5466
rect 9020 5414 9030 5466
rect 9030 5414 9076 5466
rect 8780 5412 8836 5414
rect 8860 5412 8916 5414
rect 8940 5412 8996 5414
rect 9020 5412 9076 5414
rect 8120 3834 8176 3836
rect 8200 3834 8256 3836
rect 8280 3834 8336 3836
rect 8360 3834 8416 3836
rect 8120 3782 8166 3834
rect 8166 3782 8176 3834
rect 8200 3782 8230 3834
rect 8230 3782 8242 3834
rect 8242 3782 8256 3834
rect 8280 3782 8294 3834
rect 8294 3782 8306 3834
rect 8306 3782 8336 3834
rect 8360 3782 8370 3834
rect 8370 3782 8416 3834
rect 8120 3780 8176 3782
rect 8200 3780 8256 3782
rect 8280 3780 8336 3782
rect 8360 3780 8416 3782
rect 6073 2746 6129 2748
rect 6153 2746 6209 2748
rect 6233 2746 6289 2748
rect 6313 2746 6369 2748
rect 6073 2694 6119 2746
rect 6119 2694 6129 2746
rect 6153 2694 6183 2746
rect 6183 2694 6195 2746
rect 6195 2694 6209 2746
rect 6233 2694 6247 2746
rect 6247 2694 6259 2746
rect 6259 2694 6289 2746
rect 6313 2694 6323 2746
rect 6323 2694 6369 2746
rect 6073 2692 6129 2694
rect 6153 2692 6209 2694
rect 6233 2692 6289 2694
rect 6313 2692 6369 2694
rect 8120 2746 8176 2748
rect 8200 2746 8256 2748
rect 8280 2746 8336 2748
rect 8360 2746 8416 2748
rect 8120 2694 8166 2746
rect 8166 2694 8176 2746
rect 8200 2694 8230 2746
rect 8230 2694 8242 2746
rect 8242 2694 8256 2746
rect 8280 2694 8294 2746
rect 8294 2694 8306 2746
rect 8306 2694 8336 2746
rect 8360 2694 8370 2746
rect 8370 2694 8416 2746
rect 8120 2692 8176 2694
rect 8200 2692 8256 2694
rect 8280 2692 8336 2694
rect 8360 2692 8416 2694
rect 8780 4378 8836 4380
rect 8860 4378 8916 4380
rect 8940 4378 8996 4380
rect 9020 4378 9076 4380
rect 8780 4326 8826 4378
rect 8826 4326 8836 4378
rect 8860 4326 8890 4378
rect 8890 4326 8902 4378
rect 8902 4326 8916 4378
rect 8940 4326 8954 4378
rect 8954 4326 8966 4378
rect 8966 4326 8996 4378
rect 9020 4326 9030 4378
rect 9030 4326 9076 4378
rect 8780 4324 8836 4326
rect 8860 4324 8916 4326
rect 8940 4324 8996 4326
rect 9020 4324 9076 4326
rect 8780 3290 8836 3292
rect 8860 3290 8916 3292
rect 8940 3290 8996 3292
rect 9020 3290 9076 3292
rect 8780 3238 8826 3290
rect 8826 3238 8836 3290
rect 8860 3238 8890 3290
rect 8890 3238 8902 3290
rect 8902 3238 8916 3290
rect 8940 3238 8954 3290
rect 8954 3238 8966 3290
rect 8966 3238 8996 3290
rect 9020 3238 9030 3290
rect 9030 3238 9076 3290
rect 8780 3236 8836 3238
rect 8860 3236 8916 3238
rect 8940 3236 8996 3238
rect 9020 3236 9076 3238
rect 8850 2796 8852 2816
rect 8852 2796 8904 2816
rect 8904 2796 8906 2816
rect 8850 2760 8906 2796
rect 2639 2202 2695 2204
rect 2719 2202 2775 2204
rect 2799 2202 2855 2204
rect 2879 2202 2935 2204
rect 2639 2150 2685 2202
rect 2685 2150 2695 2202
rect 2719 2150 2749 2202
rect 2749 2150 2761 2202
rect 2761 2150 2775 2202
rect 2799 2150 2813 2202
rect 2813 2150 2825 2202
rect 2825 2150 2855 2202
rect 2879 2150 2889 2202
rect 2889 2150 2935 2202
rect 2639 2148 2695 2150
rect 2719 2148 2775 2150
rect 2799 2148 2855 2150
rect 2879 2148 2935 2150
rect 4686 2202 4742 2204
rect 4766 2202 4822 2204
rect 4846 2202 4902 2204
rect 4926 2202 4982 2204
rect 4686 2150 4732 2202
rect 4732 2150 4742 2202
rect 4766 2150 4796 2202
rect 4796 2150 4808 2202
rect 4808 2150 4822 2202
rect 4846 2150 4860 2202
rect 4860 2150 4872 2202
rect 4872 2150 4902 2202
rect 4926 2150 4936 2202
rect 4936 2150 4982 2202
rect 4686 2148 4742 2150
rect 4766 2148 4822 2150
rect 4846 2148 4902 2150
rect 4926 2148 4982 2150
rect 6733 2202 6789 2204
rect 6813 2202 6869 2204
rect 6893 2202 6949 2204
rect 6973 2202 7029 2204
rect 6733 2150 6779 2202
rect 6779 2150 6789 2202
rect 6813 2150 6843 2202
rect 6843 2150 6855 2202
rect 6855 2150 6869 2202
rect 6893 2150 6907 2202
rect 6907 2150 6919 2202
rect 6919 2150 6949 2202
rect 6973 2150 6983 2202
rect 6983 2150 7029 2202
rect 6733 2148 6789 2150
rect 6813 2148 6869 2150
rect 6893 2148 6949 2150
rect 6973 2148 7029 2150
rect 8780 2202 8836 2204
rect 8860 2202 8916 2204
rect 8940 2202 8996 2204
rect 9020 2202 9076 2204
rect 8780 2150 8826 2202
rect 8826 2150 8836 2202
rect 8860 2150 8890 2202
rect 8890 2150 8902 2202
rect 8902 2150 8916 2202
rect 8940 2150 8954 2202
rect 8954 2150 8966 2202
rect 8966 2150 8996 2202
rect 9020 2150 9030 2202
rect 9030 2150 9076 2202
rect 8780 2148 8836 2150
rect 8860 2148 8916 2150
rect 8940 2148 8996 2150
rect 9020 2148 9076 2150
<< metal3 >>
rect 0 10978 800 11008
rect 933 10978 999 10981
rect 0 10976 999 10978
rect 0 10920 938 10976
rect 994 10920 999 10976
rect 0 10918 999 10920
rect 0 10888 800 10918
rect 933 10915 999 10918
rect 9213 10978 9279 10981
rect 9673 10978 10473 11008
rect 9213 10976 10473 10978
rect 9213 10920 9218 10976
rect 9274 10920 10473 10976
rect 9213 10918 10473 10920
rect 9213 10915 9279 10918
rect 9673 10888 10473 10918
rect 1969 10368 2285 10369
rect 1969 10304 1975 10368
rect 2039 10304 2055 10368
rect 2119 10304 2135 10368
rect 2199 10304 2215 10368
rect 2279 10304 2285 10368
rect 1969 10303 2285 10304
rect 4016 10368 4332 10369
rect 4016 10304 4022 10368
rect 4086 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4332 10368
rect 4016 10303 4332 10304
rect 6063 10368 6379 10369
rect 6063 10304 6069 10368
rect 6133 10304 6149 10368
rect 6213 10304 6229 10368
rect 6293 10304 6309 10368
rect 6373 10304 6379 10368
rect 6063 10303 6379 10304
rect 8110 10368 8426 10369
rect 8110 10304 8116 10368
rect 8180 10304 8196 10368
rect 8260 10304 8276 10368
rect 8340 10304 8356 10368
rect 8420 10304 8426 10368
rect 8110 10303 8426 10304
rect 2629 9824 2945 9825
rect 2629 9760 2635 9824
rect 2699 9760 2715 9824
rect 2779 9760 2795 9824
rect 2859 9760 2875 9824
rect 2939 9760 2945 9824
rect 2629 9759 2945 9760
rect 4676 9824 4992 9825
rect 4676 9760 4682 9824
rect 4746 9760 4762 9824
rect 4826 9760 4842 9824
rect 4906 9760 4922 9824
rect 4986 9760 4992 9824
rect 4676 9759 4992 9760
rect 6723 9824 7039 9825
rect 6723 9760 6729 9824
rect 6793 9760 6809 9824
rect 6873 9760 6889 9824
rect 6953 9760 6969 9824
rect 7033 9760 7039 9824
rect 6723 9759 7039 9760
rect 8770 9824 9086 9825
rect 8770 9760 8776 9824
rect 8840 9760 8856 9824
rect 8920 9760 8936 9824
rect 9000 9760 9016 9824
rect 9080 9760 9086 9824
rect 8770 9759 9086 9760
rect 1969 9280 2285 9281
rect 1969 9216 1975 9280
rect 2039 9216 2055 9280
rect 2119 9216 2135 9280
rect 2199 9216 2215 9280
rect 2279 9216 2285 9280
rect 1969 9215 2285 9216
rect 4016 9280 4332 9281
rect 4016 9216 4022 9280
rect 4086 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4332 9280
rect 4016 9215 4332 9216
rect 6063 9280 6379 9281
rect 6063 9216 6069 9280
rect 6133 9216 6149 9280
rect 6213 9216 6229 9280
rect 6293 9216 6309 9280
rect 6373 9216 6379 9280
rect 6063 9215 6379 9216
rect 8110 9280 8426 9281
rect 8110 9216 8116 9280
rect 8180 9216 8196 9280
rect 8260 9216 8276 9280
rect 8340 9216 8356 9280
rect 8420 9216 8426 9280
rect 8110 9215 8426 9216
rect 2629 8736 2945 8737
rect 2629 8672 2635 8736
rect 2699 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2875 8736
rect 2939 8672 2945 8736
rect 2629 8671 2945 8672
rect 4676 8736 4992 8737
rect 4676 8672 4682 8736
rect 4746 8672 4762 8736
rect 4826 8672 4842 8736
rect 4906 8672 4922 8736
rect 4986 8672 4992 8736
rect 4676 8671 4992 8672
rect 6723 8736 7039 8737
rect 6723 8672 6729 8736
rect 6793 8672 6809 8736
rect 6873 8672 6889 8736
rect 6953 8672 6969 8736
rect 7033 8672 7039 8736
rect 6723 8671 7039 8672
rect 8770 8736 9086 8737
rect 8770 8672 8776 8736
rect 8840 8672 8856 8736
rect 8920 8672 8936 8736
rect 9000 8672 9016 8736
rect 9080 8672 9086 8736
rect 8770 8671 9086 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 9213 8258 9279 8261
rect 9673 8258 10473 8288
rect 9213 8256 10473 8258
rect 9213 8200 9218 8256
rect 9274 8200 10473 8256
rect 9213 8198 10473 8200
rect 9213 8195 9279 8198
rect 1969 8192 2285 8193
rect 1969 8128 1975 8192
rect 2039 8128 2055 8192
rect 2119 8128 2135 8192
rect 2199 8128 2215 8192
rect 2279 8128 2285 8192
rect 1969 8127 2285 8128
rect 4016 8192 4332 8193
rect 4016 8128 4022 8192
rect 4086 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4332 8192
rect 4016 8127 4332 8128
rect 6063 8192 6379 8193
rect 6063 8128 6069 8192
rect 6133 8128 6149 8192
rect 6213 8128 6229 8192
rect 6293 8128 6309 8192
rect 6373 8128 6379 8192
rect 6063 8127 6379 8128
rect 8110 8192 8426 8193
rect 8110 8128 8116 8192
rect 8180 8128 8196 8192
rect 8260 8128 8276 8192
rect 8340 8128 8356 8192
rect 8420 8128 8426 8192
rect 9673 8168 10473 8198
rect 8110 8127 8426 8128
rect 2629 7648 2945 7649
rect 2629 7584 2635 7648
rect 2699 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2875 7648
rect 2939 7584 2945 7648
rect 2629 7583 2945 7584
rect 4676 7648 4992 7649
rect 4676 7584 4682 7648
rect 4746 7584 4762 7648
rect 4826 7584 4842 7648
rect 4906 7584 4922 7648
rect 4986 7584 4992 7648
rect 4676 7583 4992 7584
rect 6723 7648 7039 7649
rect 6723 7584 6729 7648
rect 6793 7584 6809 7648
rect 6873 7584 6889 7648
rect 6953 7584 6969 7648
rect 7033 7584 7039 7648
rect 6723 7583 7039 7584
rect 8770 7648 9086 7649
rect 8770 7584 8776 7648
rect 8840 7584 8856 7648
rect 8920 7584 8936 7648
rect 9000 7584 9016 7648
rect 9080 7584 9086 7648
rect 8770 7583 9086 7584
rect 1969 7104 2285 7105
rect 1969 7040 1975 7104
rect 2039 7040 2055 7104
rect 2119 7040 2135 7104
rect 2199 7040 2215 7104
rect 2279 7040 2285 7104
rect 1969 7039 2285 7040
rect 4016 7104 4332 7105
rect 4016 7040 4022 7104
rect 4086 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4332 7104
rect 4016 7039 4332 7040
rect 6063 7104 6379 7105
rect 6063 7040 6069 7104
rect 6133 7040 6149 7104
rect 6213 7040 6229 7104
rect 6293 7040 6309 7104
rect 6373 7040 6379 7104
rect 6063 7039 6379 7040
rect 8110 7104 8426 7105
rect 8110 7040 8116 7104
rect 8180 7040 8196 7104
rect 8260 7040 8276 7104
rect 8340 7040 8356 7104
rect 8420 7040 8426 7104
rect 8110 7039 8426 7040
rect 2629 6560 2945 6561
rect 2629 6496 2635 6560
rect 2699 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2875 6560
rect 2939 6496 2945 6560
rect 2629 6495 2945 6496
rect 4676 6560 4992 6561
rect 4676 6496 4682 6560
rect 4746 6496 4762 6560
rect 4826 6496 4842 6560
rect 4906 6496 4922 6560
rect 4986 6496 4992 6560
rect 4676 6495 4992 6496
rect 6723 6560 7039 6561
rect 6723 6496 6729 6560
rect 6793 6496 6809 6560
rect 6873 6496 6889 6560
rect 6953 6496 6969 6560
rect 7033 6496 7039 6560
rect 6723 6495 7039 6496
rect 8770 6560 9086 6561
rect 8770 6496 8776 6560
rect 8840 6496 8856 6560
rect 8920 6496 8936 6560
rect 9000 6496 9016 6560
rect 9080 6496 9086 6560
rect 8770 6495 9086 6496
rect 1969 6016 2285 6017
rect 1969 5952 1975 6016
rect 2039 5952 2055 6016
rect 2119 5952 2135 6016
rect 2199 5952 2215 6016
rect 2279 5952 2285 6016
rect 1969 5951 2285 5952
rect 4016 6016 4332 6017
rect 4016 5952 4022 6016
rect 4086 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4332 6016
rect 4016 5951 4332 5952
rect 6063 6016 6379 6017
rect 6063 5952 6069 6016
rect 6133 5952 6149 6016
rect 6213 5952 6229 6016
rect 6293 5952 6309 6016
rect 6373 5952 6379 6016
rect 6063 5951 6379 5952
rect 8110 6016 8426 6017
rect 8110 5952 8116 6016
rect 8180 5952 8196 6016
rect 8260 5952 8276 6016
rect 8340 5952 8356 6016
rect 8420 5952 8426 6016
rect 8110 5951 8426 5952
rect 4153 5810 4219 5813
rect 5441 5810 5507 5813
rect 4153 5808 5507 5810
rect 4153 5752 4158 5808
rect 4214 5752 5446 5808
rect 5502 5752 5507 5808
rect 4153 5750 5507 5752
rect 4153 5747 4219 5750
rect 5441 5747 5507 5750
rect 4337 5674 4403 5677
rect 6545 5674 6611 5677
rect 4337 5672 6611 5674
rect 4337 5616 4342 5672
rect 4398 5616 6550 5672
rect 6606 5616 6611 5672
rect 4337 5614 6611 5616
rect 4337 5611 4403 5614
rect 6545 5611 6611 5614
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 9305 5538 9371 5541
rect 9673 5538 10473 5568
rect 9305 5536 10473 5538
rect 9305 5480 9310 5536
rect 9366 5480 10473 5536
rect 9305 5478 10473 5480
rect 9305 5475 9371 5478
rect 2629 5472 2945 5473
rect 2629 5408 2635 5472
rect 2699 5408 2715 5472
rect 2779 5408 2795 5472
rect 2859 5408 2875 5472
rect 2939 5408 2945 5472
rect 2629 5407 2945 5408
rect 4676 5472 4992 5473
rect 4676 5408 4682 5472
rect 4746 5408 4762 5472
rect 4826 5408 4842 5472
rect 4906 5408 4922 5472
rect 4986 5408 4992 5472
rect 4676 5407 4992 5408
rect 6723 5472 7039 5473
rect 6723 5408 6729 5472
rect 6793 5408 6809 5472
rect 6873 5408 6889 5472
rect 6953 5408 6969 5472
rect 7033 5408 7039 5472
rect 6723 5407 7039 5408
rect 8770 5472 9086 5473
rect 8770 5408 8776 5472
rect 8840 5408 8856 5472
rect 8920 5408 8936 5472
rect 9000 5408 9016 5472
rect 9080 5408 9086 5472
rect 9673 5448 10473 5478
rect 8770 5407 9086 5408
rect 4889 5266 4955 5269
rect 7557 5266 7623 5269
rect 4889 5264 7623 5266
rect 4889 5208 4894 5264
rect 4950 5208 7562 5264
rect 7618 5208 7623 5264
rect 4889 5206 7623 5208
rect 4889 5203 4955 5206
rect 7557 5203 7623 5206
rect 1969 4928 2285 4929
rect 1969 4864 1975 4928
rect 2039 4864 2055 4928
rect 2119 4864 2135 4928
rect 2199 4864 2215 4928
rect 2279 4864 2285 4928
rect 1969 4863 2285 4864
rect 4016 4928 4332 4929
rect 4016 4864 4022 4928
rect 4086 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4332 4928
rect 4016 4863 4332 4864
rect 6063 4928 6379 4929
rect 6063 4864 6069 4928
rect 6133 4864 6149 4928
rect 6213 4864 6229 4928
rect 6293 4864 6309 4928
rect 6373 4864 6379 4928
rect 6063 4863 6379 4864
rect 8110 4928 8426 4929
rect 8110 4864 8116 4928
rect 8180 4864 8196 4928
rect 8260 4864 8276 4928
rect 8340 4864 8356 4928
rect 8420 4864 8426 4928
rect 8110 4863 8426 4864
rect 5165 4722 5231 4725
rect 5809 4722 5875 4725
rect 5165 4720 5875 4722
rect 5165 4664 5170 4720
rect 5226 4664 5814 4720
rect 5870 4664 5875 4720
rect 5165 4662 5875 4664
rect 5165 4659 5231 4662
rect 5809 4659 5875 4662
rect 2629 4384 2945 4385
rect 2629 4320 2635 4384
rect 2699 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2875 4384
rect 2939 4320 2945 4384
rect 2629 4319 2945 4320
rect 4676 4384 4992 4385
rect 4676 4320 4682 4384
rect 4746 4320 4762 4384
rect 4826 4320 4842 4384
rect 4906 4320 4922 4384
rect 4986 4320 4992 4384
rect 4676 4319 4992 4320
rect 6723 4384 7039 4385
rect 6723 4320 6729 4384
rect 6793 4320 6809 4384
rect 6873 4320 6889 4384
rect 6953 4320 6969 4384
rect 7033 4320 7039 4384
rect 6723 4319 7039 4320
rect 8770 4384 9086 4385
rect 8770 4320 8776 4384
rect 8840 4320 8856 4384
rect 8920 4320 8936 4384
rect 9000 4320 9016 4384
rect 9080 4320 9086 4384
rect 8770 4319 9086 4320
rect 1969 3840 2285 3841
rect 1969 3776 1975 3840
rect 2039 3776 2055 3840
rect 2119 3776 2135 3840
rect 2199 3776 2215 3840
rect 2279 3776 2285 3840
rect 1969 3775 2285 3776
rect 4016 3840 4332 3841
rect 4016 3776 4022 3840
rect 4086 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4332 3840
rect 4016 3775 4332 3776
rect 6063 3840 6379 3841
rect 6063 3776 6069 3840
rect 6133 3776 6149 3840
rect 6213 3776 6229 3840
rect 6293 3776 6309 3840
rect 6373 3776 6379 3840
rect 6063 3775 6379 3776
rect 8110 3840 8426 3841
rect 8110 3776 8116 3840
rect 8180 3776 8196 3840
rect 8260 3776 8276 3840
rect 8340 3776 8356 3840
rect 8420 3776 8426 3840
rect 8110 3775 8426 3776
rect 2629 3296 2945 3297
rect 2629 3232 2635 3296
rect 2699 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2875 3296
rect 2939 3232 2945 3296
rect 2629 3231 2945 3232
rect 4676 3296 4992 3297
rect 4676 3232 4682 3296
rect 4746 3232 4762 3296
rect 4826 3232 4842 3296
rect 4906 3232 4922 3296
rect 4986 3232 4992 3296
rect 4676 3231 4992 3232
rect 6723 3296 7039 3297
rect 6723 3232 6729 3296
rect 6793 3232 6809 3296
rect 6873 3232 6889 3296
rect 6953 3232 6969 3296
rect 7033 3232 7039 3296
rect 6723 3231 7039 3232
rect 8770 3296 9086 3297
rect 8770 3232 8776 3296
rect 8840 3232 8856 3296
rect 8920 3232 8936 3296
rect 9000 3232 9016 3296
rect 9080 3232 9086 3296
rect 8770 3231 9086 3232
rect 2497 2954 2563 2957
rect 5257 2954 5323 2957
rect 2497 2952 5323 2954
rect 2497 2896 2502 2952
rect 2558 2896 5262 2952
rect 5318 2896 5323 2952
rect 2497 2894 5323 2896
rect 2497 2891 2563 2894
rect 5257 2891 5323 2894
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 8845 2818 8911 2821
rect 9673 2818 10473 2848
rect 8845 2816 10473 2818
rect 8845 2760 8850 2816
rect 8906 2760 10473 2816
rect 8845 2758 10473 2760
rect 8845 2755 8911 2758
rect 1969 2752 2285 2753
rect 1969 2688 1975 2752
rect 2039 2688 2055 2752
rect 2119 2688 2135 2752
rect 2199 2688 2215 2752
rect 2279 2688 2285 2752
rect 1969 2687 2285 2688
rect 4016 2752 4332 2753
rect 4016 2688 4022 2752
rect 4086 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4332 2752
rect 4016 2687 4332 2688
rect 6063 2752 6379 2753
rect 6063 2688 6069 2752
rect 6133 2688 6149 2752
rect 6213 2688 6229 2752
rect 6293 2688 6309 2752
rect 6373 2688 6379 2752
rect 6063 2687 6379 2688
rect 8110 2752 8426 2753
rect 8110 2688 8116 2752
rect 8180 2688 8196 2752
rect 8260 2688 8276 2752
rect 8340 2688 8356 2752
rect 8420 2688 8426 2752
rect 9673 2728 10473 2758
rect 8110 2687 8426 2688
rect 2629 2208 2945 2209
rect 2629 2144 2635 2208
rect 2699 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2875 2208
rect 2939 2144 2945 2208
rect 2629 2143 2945 2144
rect 4676 2208 4992 2209
rect 4676 2144 4682 2208
rect 4746 2144 4762 2208
rect 4826 2144 4842 2208
rect 4906 2144 4922 2208
rect 4986 2144 4992 2208
rect 4676 2143 4992 2144
rect 6723 2208 7039 2209
rect 6723 2144 6729 2208
rect 6793 2144 6809 2208
rect 6873 2144 6889 2208
rect 6953 2144 6969 2208
rect 7033 2144 7039 2208
rect 6723 2143 7039 2144
rect 8770 2208 9086 2209
rect 8770 2144 8776 2208
rect 8840 2144 8856 2208
rect 8920 2144 8936 2208
rect 9000 2144 9016 2208
rect 9080 2144 9086 2208
rect 8770 2143 9086 2144
<< via3 >>
rect 1975 10364 2039 10368
rect 1975 10308 1979 10364
rect 1979 10308 2035 10364
rect 2035 10308 2039 10364
rect 1975 10304 2039 10308
rect 2055 10364 2119 10368
rect 2055 10308 2059 10364
rect 2059 10308 2115 10364
rect 2115 10308 2119 10364
rect 2055 10304 2119 10308
rect 2135 10364 2199 10368
rect 2135 10308 2139 10364
rect 2139 10308 2195 10364
rect 2195 10308 2199 10364
rect 2135 10304 2199 10308
rect 2215 10364 2279 10368
rect 2215 10308 2219 10364
rect 2219 10308 2275 10364
rect 2275 10308 2279 10364
rect 2215 10304 2279 10308
rect 4022 10364 4086 10368
rect 4022 10308 4026 10364
rect 4026 10308 4082 10364
rect 4082 10308 4086 10364
rect 4022 10304 4086 10308
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 6069 10364 6133 10368
rect 6069 10308 6073 10364
rect 6073 10308 6129 10364
rect 6129 10308 6133 10364
rect 6069 10304 6133 10308
rect 6149 10364 6213 10368
rect 6149 10308 6153 10364
rect 6153 10308 6209 10364
rect 6209 10308 6213 10364
rect 6149 10304 6213 10308
rect 6229 10364 6293 10368
rect 6229 10308 6233 10364
rect 6233 10308 6289 10364
rect 6289 10308 6293 10364
rect 6229 10304 6293 10308
rect 6309 10364 6373 10368
rect 6309 10308 6313 10364
rect 6313 10308 6369 10364
rect 6369 10308 6373 10364
rect 6309 10304 6373 10308
rect 8116 10364 8180 10368
rect 8116 10308 8120 10364
rect 8120 10308 8176 10364
rect 8176 10308 8180 10364
rect 8116 10304 8180 10308
rect 8196 10364 8260 10368
rect 8196 10308 8200 10364
rect 8200 10308 8256 10364
rect 8256 10308 8260 10364
rect 8196 10304 8260 10308
rect 8276 10364 8340 10368
rect 8276 10308 8280 10364
rect 8280 10308 8336 10364
rect 8336 10308 8340 10364
rect 8276 10304 8340 10308
rect 8356 10364 8420 10368
rect 8356 10308 8360 10364
rect 8360 10308 8416 10364
rect 8416 10308 8420 10364
rect 8356 10304 8420 10308
rect 2635 9820 2699 9824
rect 2635 9764 2639 9820
rect 2639 9764 2695 9820
rect 2695 9764 2699 9820
rect 2635 9760 2699 9764
rect 2715 9820 2779 9824
rect 2715 9764 2719 9820
rect 2719 9764 2775 9820
rect 2775 9764 2779 9820
rect 2715 9760 2779 9764
rect 2795 9820 2859 9824
rect 2795 9764 2799 9820
rect 2799 9764 2855 9820
rect 2855 9764 2859 9820
rect 2795 9760 2859 9764
rect 2875 9820 2939 9824
rect 2875 9764 2879 9820
rect 2879 9764 2935 9820
rect 2935 9764 2939 9820
rect 2875 9760 2939 9764
rect 4682 9820 4746 9824
rect 4682 9764 4686 9820
rect 4686 9764 4742 9820
rect 4742 9764 4746 9820
rect 4682 9760 4746 9764
rect 4762 9820 4826 9824
rect 4762 9764 4766 9820
rect 4766 9764 4822 9820
rect 4822 9764 4826 9820
rect 4762 9760 4826 9764
rect 4842 9820 4906 9824
rect 4842 9764 4846 9820
rect 4846 9764 4902 9820
rect 4902 9764 4906 9820
rect 4842 9760 4906 9764
rect 4922 9820 4986 9824
rect 4922 9764 4926 9820
rect 4926 9764 4982 9820
rect 4982 9764 4986 9820
rect 4922 9760 4986 9764
rect 6729 9820 6793 9824
rect 6729 9764 6733 9820
rect 6733 9764 6789 9820
rect 6789 9764 6793 9820
rect 6729 9760 6793 9764
rect 6809 9820 6873 9824
rect 6809 9764 6813 9820
rect 6813 9764 6869 9820
rect 6869 9764 6873 9820
rect 6809 9760 6873 9764
rect 6889 9820 6953 9824
rect 6889 9764 6893 9820
rect 6893 9764 6949 9820
rect 6949 9764 6953 9820
rect 6889 9760 6953 9764
rect 6969 9820 7033 9824
rect 6969 9764 6973 9820
rect 6973 9764 7029 9820
rect 7029 9764 7033 9820
rect 6969 9760 7033 9764
rect 8776 9820 8840 9824
rect 8776 9764 8780 9820
rect 8780 9764 8836 9820
rect 8836 9764 8840 9820
rect 8776 9760 8840 9764
rect 8856 9820 8920 9824
rect 8856 9764 8860 9820
rect 8860 9764 8916 9820
rect 8916 9764 8920 9820
rect 8856 9760 8920 9764
rect 8936 9820 9000 9824
rect 8936 9764 8940 9820
rect 8940 9764 8996 9820
rect 8996 9764 9000 9820
rect 8936 9760 9000 9764
rect 9016 9820 9080 9824
rect 9016 9764 9020 9820
rect 9020 9764 9076 9820
rect 9076 9764 9080 9820
rect 9016 9760 9080 9764
rect 1975 9276 2039 9280
rect 1975 9220 1979 9276
rect 1979 9220 2035 9276
rect 2035 9220 2039 9276
rect 1975 9216 2039 9220
rect 2055 9276 2119 9280
rect 2055 9220 2059 9276
rect 2059 9220 2115 9276
rect 2115 9220 2119 9276
rect 2055 9216 2119 9220
rect 2135 9276 2199 9280
rect 2135 9220 2139 9276
rect 2139 9220 2195 9276
rect 2195 9220 2199 9276
rect 2135 9216 2199 9220
rect 2215 9276 2279 9280
rect 2215 9220 2219 9276
rect 2219 9220 2275 9276
rect 2275 9220 2279 9276
rect 2215 9216 2279 9220
rect 4022 9276 4086 9280
rect 4022 9220 4026 9276
rect 4026 9220 4082 9276
rect 4082 9220 4086 9276
rect 4022 9216 4086 9220
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 6069 9276 6133 9280
rect 6069 9220 6073 9276
rect 6073 9220 6129 9276
rect 6129 9220 6133 9276
rect 6069 9216 6133 9220
rect 6149 9276 6213 9280
rect 6149 9220 6153 9276
rect 6153 9220 6209 9276
rect 6209 9220 6213 9276
rect 6149 9216 6213 9220
rect 6229 9276 6293 9280
rect 6229 9220 6233 9276
rect 6233 9220 6289 9276
rect 6289 9220 6293 9276
rect 6229 9216 6293 9220
rect 6309 9276 6373 9280
rect 6309 9220 6313 9276
rect 6313 9220 6369 9276
rect 6369 9220 6373 9276
rect 6309 9216 6373 9220
rect 8116 9276 8180 9280
rect 8116 9220 8120 9276
rect 8120 9220 8176 9276
rect 8176 9220 8180 9276
rect 8116 9216 8180 9220
rect 8196 9276 8260 9280
rect 8196 9220 8200 9276
rect 8200 9220 8256 9276
rect 8256 9220 8260 9276
rect 8196 9216 8260 9220
rect 8276 9276 8340 9280
rect 8276 9220 8280 9276
rect 8280 9220 8336 9276
rect 8336 9220 8340 9276
rect 8276 9216 8340 9220
rect 8356 9276 8420 9280
rect 8356 9220 8360 9276
rect 8360 9220 8416 9276
rect 8416 9220 8420 9276
rect 8356 9216 8420 9220
rect 2635 8732 2699 8736
rect 2635 8676 2639 8732
rect 2639 8676 2695 8732
rect 2695 8676 2699 8732
rect 2635 8672 2699 8676
rect 2715 8732 2779 8736
rect 2715 8676 2719 8732
rect 2719 8676 2775 8732
rect 2775 8676 2779 8732
rect 2715 8672 2779 8676
rect 2795 8732 2859 8736
rect 2795 8676 2799 8732
rect 2799 8676 2855 8732
rect 2855 8676 2859 8732
rect 2795 8672 2859 8676
rect 2875 8732 2939 8736
rect 2875 8676 2879 8732
rect 2879 8676 2935 8732
rect 2935 8676 2939 8732
rect 2875 8672 2939 8676
rect 4682 8732 4746 8736
rect 4682 8676 4686 8732
rect 4686 8676 4742 8732
rect 4742 8676 4746 8732
rect 4682 8672 4746 8676
rect 4762 8732 4826 8736
rect 4762 8676 4766 8732
rect 4766 8676 4822 8732
rect 4822 8676 4826 8732
rect 4762 8672 4826 8676
rect 4842 8732 4906 8736
rect 4842 8676 4846 8732
rect 4846 8676 4902 8732
rect 4902 8676 4906 8732
rect 4842 8672 4906 8676
rect 4922 8732 4986 8736
rect 4922 8676 4926 8732
rect 4926 8676 4982 8732
rect 4982 8676 4986 8732
rect 4922 8672 4986 8676
rect 6729 8732 6793 8736
rect 6729 8676 6733 8732
rect 6733 8676 6789 8732
rect 6789 8676 6793 8732
rect 6729 8672 6793 8676
rect 6809 8732 6873 8736
rect 6809 8676 6813 8732
rect 6813 8676 6869 8732
rect 6869 8676 6873 8732
rect 6809 8672 6873 8676
rect 6889 8732 6953 8736
rect 6889 8676 6893 8732
rect 6893 8676 6949 8732
rect 6949 8676 6953 8732
rect 6889 8672 6953 8676
rect 6969 8732 7033 8736
rect 6969 8676 6973 8732
rect 6973 8676 7029 8732
rect 7029 8676 7033 8732
rect 6969 8672 7033 8676
rect 8776 8732 8840 8736
rect 8776 8676 8780 8732
rect 8780 8676 8836 8732
rect 8836 8676 8840 8732
rect 8776 8672 8840 8676
rect 8856 8732 8920 8736
rect 8856 8676 8860 8732
rect 8860 8676 8916 8732
rect 8916 8676 8920 8732
rect 8856 8672 8920 8676
rect 8936 8732 9000 8736
rect 8936 8676 8940 8732
rect 8940 8676 8996 8732
rect 8996 8676 9000 8732
rect 8936 8672 9000 8676
rect 9016 8732 9080 8736
rect 9016 8676 9020 8732
rect 9020 8676 9076 8732
rect 9076 8676 9080 8732
rect 9016 8672 9080 8676
rect 1975 8188 2039 8192
rect 1975 8132 1979 8188
rect 1979 8132 2035 8188
rect 2035 8132 2039 8188
rect 1975 8128 2039 8132
rect 2055 8188 2119 8192
rect 2055 8132 2059 8188
rect 2059 8132 2115 8188
rect 2115 8132 2119 8188
rect 2055 8128 2119 8132
rect 2135 8188 2199 8192
rect 2135 8132 2139 8188
rect 2139 8132 2195 8188
rect 2195 8132 2199 8188
rect 2135 8128 2199 8132
rect 2215 8188 2279 8192
rect 2215 8132 2219 8188
rect 2219 8132 2275 8188
rect 2275 8132 2279 8188
rect 2215 8128 2279 8132
rect 4022 8188 4086 8192
rect 4022 8132 4026 8188
rect 4026 8132 4082 8188
rect 4082 8132 4086 8188
rect 4022 8128 4086 8132
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 6069 8188 6133 8192
rect 6069 8132 6073 8188
rect 6073 8132 6129 8188
rect 6129 8132 6133 8188
rect 6069 8128 6133 8132
rect 6149 8188 6213 8192
rect 6149 8132 6153 8188
rect 6153 8132 6209 8188
rect 6209 8132 6213 8188
rect 6149 8128 6213 8132
rect 6229 8188 6293 8192
rect 6229 8132 6233 8188
rect 6233 8132 6289 8188
rect 6289 8132 6293 8188
rect 6229 8128 6293 8132
rect 6309 8188 6373 8192
rect 6309 8132 6313 8188
rect 6313 8132 6369 8188
rect 6369 8132 6373 8188
rect 6309 8128 6373 8132
rect 8116 8188 8180 8192
rect 8116 8132 8120 8188
rect 8120 8132 8176 8188
rect 8176 8132 8180 8188
rect 8116 8128 8180 8132
rect 8196 8188 8260 8192
rect 8196 8132 8200 8188
rect 8200 8132 8256 8188
rect 8256 8132 8260 8188
rect 8196 8128 8260 8132
rect 8276 8188 8340 8192
rect 8276 8132 8280 8188
rect 8280 8132 8336 8188
rect 8336 8132 8340 8188
rect 8276 8128 8340 8132
rect 8356 8188 8420 8192
rect 8356 8132 8360 8188
rect 8360 8132 8416 8188
rect 8416 8132 8420 8188
rect 8356 8128 8420 8132
rect 2635 7644 2699 7648
rect 2635 7588 2639 7644
rect 2639 7588 2695 7644
rect 2695 7588 2699 7644
rect 2635 7584 2699 7588
rect 2715 7644 2779 7648
rect 2715 7588 2719 7644
rect 2719 7588 2775 7644
rect 2775 7588 2779 7644
rect 2715 7584 2779 7588
rect 2795 7644 2859 7648
rect 2795 7588 2799 7644
rect 2799 7588 2855 7644
rect 2855 7588 2859 7644
rect 2795 7584 2859 7588
rect 2875 7644 2939 7648
rect 2875 7588 2879 7644
rect 2879 7588 2935 7644
rect 2935 7588 2939 7644
rect 2875 7584 2939 7588
rect 4682 7644 4746 7648
rect 4682 7588 4686 7644
rect 4686 7588 4742 7644
rect 4742 7588 4746 7644
rect 4682 7584 4746 7588
rect 4762 7644 4826 7648
rect 4762 7588 4766 7644
rect 4766 7588 4822 7644
rect 4822 7588 4826 7644
rect 4762 7584 4826 7588
rect 4842 7644 4906 7648
rect 4842 7588 4846 7644
rect 4846 7588 4902 7644
rect 4902 7588 4906 7644
rect 4842 7584 4906 7588
rect 4922 7644 4986 7648
rect 4922 7588 4926 7644
rect 4926 7588 4982 7644
rect 4982 7588 4986 7644
rect 4922 7584 4986 7588
rect 6729 7644 6793 7648
rect 6729 7588 6733 7644
rect 6733 7588 6789 7644
rect 6789 7588 6793 7644
rect 6729 7584 6793 7588
rect 6809 7644 6873 7648
rect 6809 7588 6813 7644
rect 6813 7588 6869 7644
rect 6869 7588 6873 7644
rect 6809 7584 6873 7588
rect 6889 7644 6953 7648
rect 6889 7588 6893 7644
rect 6893 7588 6949 7644
rect 6949 7588 6953 7644
rect 6889 7584 6953 7588
rect 6969 7644 7033 7648
rect 6969 7588 6973 7644
rect 6973 7588 7029 7644
rect 7029 7588 7033 7644
rect 6969 7584 7033 7588
rect 8776 7644 8840 7648
rect 8776 7588 8780 7644
rect 8780 7588 8836 7644
rect 8836 7588 8840 7644
rect 8776 7584 8840 7588
rect 8856 7644 8920 7648
rect 8856 7588 8860 7644
rect 8860 7588 8916 7644
rect 8916 7588 8920 7644
rect 8856 7584 8920 7588
rect 8936 7644 9000 7648
rect 8936 7588 8940 7644
rect 8940 7588 8996 7644
rect 8996 7588 9000 7644
rect 8936 7584 9000 7588
rect 9016 7644 9080 7648
rect 9016 7588 9020 7644
rect 9020 7588 9076 7644
rect 9076 7588 9080 7644
rect 9016 7584 9080 7588
rect 1975 7100 2039 7104
rect 1975 7044 1979 7100
rect 1979 7044 2035 7100
rect 2035 7044 2039 7100
rect 1975 7040 2039 7044
rect 2055 7100 2119 7104
rect 2055 7044 2059 7100
rect 2059 7044 2115 7100
rect 2115 7044 2119 7100
rect 2055 7040 2119 7044
rect 2135 7100 2199 7104
rect 2135 7044 2139 7100
rect 2139 7044 2195 7100
rect 2195 7044 2199 7100
rect 2135 7040 2199 7044
rect 2215 7100 2279 7104
rect 2215 7044 2219 7100
rect 2219 7044 2275 7100
rect 2275 7044 2279 7100
rect 2215 7040 2279 7044
rect 4022 7100 4086 7104
rect 4022 7044 4026 7100
rect 4026 7044 4082 7100
rect 4082 7044 4086 7100
rect 4022 7040 4086 7044
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 6069 7100 6133 7104
rect 6069 7044 6073 7100
rect 6073 7044 6129 7100
rect 6129 7044 6133 7100
rect 6069 7040 6133 7044
rect 6149 7100 6213 7104
rect 6149 7044 6153 7100
rect 6153 7044 6209 7100
rect 6209 7044 6213 7100
rect 6149 7040 6213 7044
rect 6229 7100 6293 7104
rect 6229 7044 6233 7100
rect 6233 7044 6289 7100
rect 6289 7044 6293 7100
rect 6229 7040 6293 7044
rect 6309 7100 6373 7104
rect 6309 7044 6313 7100
rect 6313 7044 6369 7100
rect 6369 7044 6373 7100
rect 6309 7040 6373 7044
rect 8116 7100 8180 7104
rect 8116 7044 8120 7100
rect 8120 7044 8176 7100
rect 8176 7044 8180 7100
rect 8116 7040 8180 7044
rect 8196 7100 8260 7104
rect 8196 7044 8200 7100
rect 8200 7044 8256 7100
rect 8256 7044 8260 7100
rect 8196 7040 8260 7044
rect 8276 7100 8340 7104
rect 8276 7044 8280 7100
rect 8280 7044 8336 7100
rect 8336 7044 8340 7100
rect 8276 7040 8340 7044
rect 8356 7100 8420 7104
rect 8356 7044 8360 7100
rect 8360 7044 8416 7100
rect 8416 7044 8420 7100
rect 8356 7040 8420 7044
rect 2635 6556 2699 6560
rect 2635 6500 2639 6556
rect 2639 6500 2695 6556
rect 2695 6500 2699 6556
rect 2635 6496 2699 6500
rect 2715 6556 2779 6560
rect 2715 6500 2719 6556
rect 2719 6500 2775 6556
rect 2775 6500 2779 6556
rect 2715 6496 2779 6500
rect 2795 6556 2859 6560
rect 2795 6500 2799 6556
rect 2799 6500 2855 6556
rect 2855 6500 2859 6556
rect 2795 6496 2859 6500
rect 2875 6556 2939 6560
rect 2875 6500 2879 6556
rect 2879 6500 2935 6556
rect 2935 6500 2939 6556
rect 2875 6496 2939 6500
rect 4682 6556 4746 6560
rect 4682 6500 4686 6556
rect 4686 6500 4742 6556
rect 4742 6500 4746 6556
rect 4682 6496 4746 6500
rect 4762 6556 4826 6560
rect 4762 6500 4766 6556
rect 4766 6500 4822 6556
rect 4822 6500 4826 6556
rect 4762 6496 4826 6500
rect 4842 6556 4906 6560
rect 4842 6500 4846 6556
rect 4846 6500 4902 6556
rect 4902 6500 4906 6556
rect 4842 6496 4906 6500
rect 4922 6556 4986 6560
rect 4922 6500 4926 6556
rect 4926 6500 4982 6556
rect 4982 6500 4986 6556
rect 4922 6496 4986 6500
rect 6729 6556 6793 6560
rect 6729 6500 6733 6556
rect 6733 6500 6789 6556
rect 6789 6500 6793 6556
rect 6729 6496 6793 6500
rect 6809 6556 6873 6560
rect 6809 6500 6813 6556
rect 6813 6500 6869 6556
rect 6869 6500 6873 6556
rect 6809 6496 6873 6500
rect 6889 6556 6953 6560
rect 6889 6500 6893 6556
rect 6893 6500 6949 6556
rect 6949 6500 6953 6556
rect 6889 6496 6953 6500
rect 6969 6556 7033 6560
rect 6969 6500 6973 6556
rect 6973 6500 7029 6556
rect 7029 6500 7033 6556
rect 6969 6496 7033 6500
rect 8776 6556 8840 6560
rect 8776 6500 8780 6556
rect 8780 6500 8836 6556
rect 8836 6500 8840 6556
rect 8776 6496 8840 6500
rect 8856 6556 8920 6560
rect 8856 6500 8860 6556
rect 8860 6500 8916 6556
rect 8916 6500 8920 6556
rect 8856 6496 8920 6500
rect 8936 6556 9000 6560
rect 8936 6500 8940 6556
rect 8940 6500 8996 6556
rect 8996 6500 9000 6556
rect 8936 6496 9000 6500
rect 9016 6556 9080 6560
rect 9016 6500 9020 6556
rect 9020 6500 9076 6556
rect 9076 6500 9080 6556
rect 9016 6496 9080 6500
rect 1975 6012 2039 6016
rect 1975 5956 1979 6012
rect 1979 5956 2035 6012
rect 2035 5956 2039 6012
rect 1975 5952 2039 5956
rect 2055 6012 2119 6016
rect 2055 5956 2059 6012
rect 2059 5956 2115 6012
rect 2115 5956 2119 6012
rect 2055 5952 2119 5956
rect 2135 6012 2199 6016
rect 2135 5956 2139 6012
rect 2139 5956 2195 6012
rect 2195 5956 2199 6012
rect 2135 5952 2199 5956
rect 2215 6012 2279 6016
rect 2215 5956 2219 6012
rect 2219 5956 2275 6012
rect 2275 5956 2279 6012
rect 2215 5952 2279 5956
rect 4022 6012 4086 6016
rect 4022 5956 4026 6012
rect 4026 5956 4082 6012
rect 4082 5956 4086 6012
rect 4022 5952 4086 5956
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 6069 6012 6133 6016
rect 6069 5956 6073 6012
rect 6073 5956 6129 6012
rect 6129 5956 6133 6012
rect 6069 5952 6133 5956
rect 6149 6012 6213 6016
rect 6149 5956 6153 6012
rect 6153 5956 6209 6012
rect 6209 5956 6213 6012
rect 6149 5952 6213 5956
rect 6229 6012 6293 6016
rect 6229 5956 6233 6012
rect 6233 5956 6289 6012
rect 6289 5956 6293 6012
rect 6229 5952 6293 5956
rect 6309 6012 6373 6016
rect 6309 5956 6313 6012
rect 6313 5956 6369 6012
rect 6369 5956 6373 6012
rect 6309 5952 6373 5956
rect 8116 6012 8180 6016
rect 8116 5956 8120 6012
rect 8120 5956 8176 6012
rect 8176 5956 8180 6012
rect 8116 5952 8180 5956
rect 8196 6012 8260 6016
rect 8196 5956 8200 6012
rect 8200 5956 8256 6012
rect 8256 5956 8260 6012
rect 8196 5952 8260 5956
rect 8276 6012 8340 6016
rect 8276 5956 8280 6012
rect 8280 5956 8336 6012
rect 8336 5956 8340 6012
rect 8276 5952 8340 5956
rect 8356 6012 8420 6016
rect 8356 5956 8360 6012
rect 8360 5956 8416 6012
rect 8416 5956 8420 6012
rect 8356 5952 8420 5956
rect 2635 5468 2699 5472
rect 2635 5412 2639 5468
rect 2639 5412 2695 5468
rect 2695 5412 2699 5468
rect 2635 5408 2699 5412
rect 2715 5468 2779 5472
rect 2715 5412 2719 5468
rect 2719 5412 2775 5468
rect 2775 5412 2779 5468
rect 2715 5408 2779 5412
rect 2795 5468 2859 5472
rect 2795 5412 2799 5468
rect 2799 5412 2855 5468
rect 2855 5412 2859 5468
rect 2795 5408 2859 5412
rect 2875 5468 2939 5472
rect 2875 5412 2879 5468
rect 2879 5412 2935 5468
rect 2935 5412 2939 5468
rect 2875 5408 2939 5412
rect 4682 5468 4746 5472
rect 4682 5412 4686 5468
rect 4686 5412 4742 5468
rect 4742 5412 4746 5468
rect 4682 5408 4746 5412
rect 4762 5468 4826 5472
rect 4762 5412 4766 5468
rect 4766 5412 4822 5468
rect 4822 5412 4826 5468
rect 4762 5408 4826 5412
rect 4842 5468 4906 5472
rect 4842 5412 4846 5468
rect 4846 5412 4902 5468
rect 4902 5412 4906 5468
rect 4842 5408 4906 5412
rect 4922 5468 4986 5472
rect 4922 5412 4926 5468
rect 4926 5412 4982 5468
rect 4982 5412 4986 5468
rect 4922 5408 4986 5412
rect 6729 5468 6793 5472
rect 6729 5412 6733 5468
rect 6733 5412 6789 5468
rect 6789 5412 6793 5468
rect 6729 5408 6793 5412
rect 6809 5468 6873 5472
rect 6809 5412 6813 5468
rect 6813 5412 6869 5468
rect 6869 5412 6873 5468
rect 6809 5408 6873 5412
rect 6889 5468 6953 5472
rect 6889 5412 6893 5468
rect 6893 5412 6949 5468
rect 6949 5412 6953 5468
rect 6889 5408 6953 5412
rect 6969 5468 7033 5472
rect 6969 5412 6973 5468
rect 6973 5412 7029 5468
rect 7029 5412 7033 5468
rect 6969 5408 7033 5412
rect 8776 5468 8840 5472
rect 8776 5412 8780 5468
rect 8780 5412 8836 5468
rect 8836 5412 8840 5468
rect 8776 5408 8840 5412
rect 8856 5468 8920 5472
rect 8856 5412 8860 5468
rect 8860 5412 8916 5468
rect 8916 5412 8920 5468
rect 8856 5408 8920 5412
rect 8936 5468 9000 5472
rect 8936 5412 8940 5468
rect 8940 5412 8996 5468
rect 8996 5412 9000 5468
rect 8936 5408 9000 5412
rect 9016 5468 9080 5472
rect 9016 5412 9020 5468
rect 9020 5412 9076 5468
rect 9076 5412 9080 5468
rect 9016 5408 9080 5412
rect 1975 4924 2039 4928
rect 1975 4868 1979 4924
rect 1979 4868 2035 4924
rect 2035 4868 2039 4924
rect 1975 4864 2039 4868
rect 2055 4924 2119 4928
rect 2055 4868 2059 4924
rect 2059 4868 2115 4924
rect 2115 4868 2119 4924
rect 2055 4864 2119 4868
rect 2135 4924 2199 4928
rect 2135 4868 2139 4924
rect 2139 4868 2195 4924
rect 2195 4868 2199 4924
rect 2135 4864 2199 4868
rect 2215 4924 2279 4928
rect 2215 4868 2219 4924
rect 2219 4868 2275 4924
rect 2275 4868 2279 4924
rect 2215 4864 2279 4868
rect 4022 4924 4086 4928
rect 4022 4868 4026 4924
rect 4026 4868 4082 4924
rect 4082 4868 4086 4924
rect 4022 4864 4086 4868
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 6069 4924 6133 4928
rect 6069 4868 6073 4924
rect 6073 4868 6129 4924
rect 6129 4868 6133 4924
rect 6069 4864 6133 4868
rect 6149 4924 6213 4928
rect 6149 4868 6153 4924
rect 6153 4868 6209 4924
rect 6209 4868 6213 4924
rect 6149 4864 6213 4868
rect 6229 4924 6293 4928
rect 6229 4868 6233 4924
rect 6233 4868 6289 4924
rect 6289 4868 6293 4924
rect 6229 4864 6293 4868
rect 6309 4924 6373 4928
rect 6309 4868 6313 4924
rect 6313 4868 6369 4924
rect 6369 4868 6373 4924
rect 6309 4864 6373 4868
rect 8116 4924 8180 4928
rect 8116 4868 8120 4924
rect 8120 4868 8176 4924
rect 8176 4868 8180 4924
rect 8116 4864 8180 4868
rect 8196 4924 8260 4928
rect 8196 4868 8200 4924
rect 8200 4868 8256 4924
rect 8256 4868 8260 4924
rect 8196 4864 8260 4868
rect 8276 4924 8340 4928
rect 8276 4868 8280 4924
rect 8280 4868 8336 4924
rect 8336 4868 8340 4924
rect 8276 4864 8340 4868
rect 8356 4924 8420 4928
rect 8356 4868 8360 4924
rect 8360 4868 8416 4924
rect 8416 4868 8420 4924
rect 8356 4864 8420 4868
rect 2635 4380 2699 4384
rect 2635 4324 2639 4380
rect 2639 4324 2695 4380
rect 2695 4324 2699 4380
rect 2635 4320 2699 4324
rect 2715 4380 2779 4384
rect 2715 4324 2719 4380
rect 2719 4324 2775 4380
rect 2775 4324 2779 4380
rect 2715 4320 2779 4324
rect 2795 4380 2859 4384
rect 2795 4324 2799 4380
rect 2799 4324 2855 4380
rect 2855 4324 2859 4380
rect 2795 4320 2859 4324
rect 2875 4380 2939 4384
rect 2875 4324 2879 4380
rect 2879 4324 2935 4380
rect 2935 4324 2939 4380
rect 2875 4320 2939 4324
rect 4682 4380 4746 4384
rect 4682 4324 4686 4380
rect 4686 4324 4742 4380
rect 4742 4324 4746 4380
rect 4682 4320 4746 4324
rect 4762 4380 4826 4384
rect 4762 4324 4766 4380
rect 4766 4324 4822 4380
rect 4822 4324 4826 4380
rect 4762 4320 4826 4324
rect 4842 4380 4906 4384
rect 4842 4324 4846 4380
rect 4846 4324 4902 4380
rect 4902 4324 4906 4380
rect 4842 4320 4906 4324
rect 4922 4380 4986 4384
rect 4922 4324 4926 4380
rect 4926 4324 4982 4380
rect 4982 4324 4986 4380
rect 4922 4320 4986 4324
rect 6729 4380 6793 4384
rect 6729 4324 6733 4380
rect 6733 4324 6789 4380
rect 6789 4324 6793 4380
rect 6729 4320 6793 4324
rect 6809 4380 6873 4384
rect 6809 4324 6813 4380
rect 6813 4324 6869 4380
rect 6869 4324 6873 4380
rect 6809 4320 6873 4324
rect 6889 4380 6953 4384
rect 6889 4324 6893 4380
rect 6893 4324 6949 4380
rect 6949 4324 6953 4380
rect 6889 4320 6953 4324
rect 6969 4380 7033 4384
rect 6969 4324 6973 4380
rect 6973 4324 7029 4380
rect 7029 4324 7033 4380
rect 6969 4320 7033 4324
rect 8776 4380 8840 4384
rect 8776 4324 8780 4380
rect 8780 4324 8836 4380
rect 8836 4324 8840 4380
rect 8776 4320 8840 4324
rect 8856 4380 8920 4384
rect 8856 4324 8860 4380
rect 8860 4324 8916 4380
rect 8916 4324 8920 4380
rect 8856 4320 8920 4324
rect 8936 4380 9000 4384
rect 8936 4324 8940 4380
rect 8940 4324 8996 4380
rect 8996 4324 9000 4380
rect 8936 4320 9000 4324
rect 9016 4380 9080 4384
rect 9016 4324 9020 4380
rect 9020 4324 9076 4380
rect 9076 4324 9080 4380
rect 9016 4320 9080 4324
rect 1975 3836 2039 3840
rect 1975 3780 1979 3836
rect 1979 3780 2035 3836
rect 2035 3780 2039 3836
rect 1975 3776 2039 3780
rect 2055 3836 2119 3840
rect 2055 3780 2059 3836
rect 2059 3780 2115 3836
rect 2115 3780 2119 3836
rect 2055 3776 2119 3780
rect 2135 3836 2199 3840
rect 2135 3780 2139 3836
rect 2139 3780 2195 3836
rect 2195 3780 2199 3836
rect 2135 3776 2199 3780
rect 2215 3836 2279 3840
rect 2215 3780 2219 3836
rect 2219 3780 2275 3836
rect 2275 3780 2279 3836
rect 2215 3776 2279 3780
rect 4022 3836 4086 3840
rect 4022 3780 4026 3836
rect 4026 3780 4082 3836
rect 4082 3780 4086 3836
rect 4022 3776 4086 3780
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 6069 3836 6133 3840
rect 6069 3780 6073 3836
rect 6073 3780 6129 3836
rect 6129 3780 6133 3836
rect 6069 3776 6133 3780
rect 6149 3836 6213 3840
rect 6149 3780 6153 3836
rect 6153 3780 6209 3836
rect 6209 3780 6213 3836
rect 6149 3776 6213 3780
rect 6229 3836 6293 3840
rect 6229 3780 6233 3836
rect 6233 3780 6289 3836
rect 6289 3780 6293 3836
rect 6229 3776 6293 3780
rect 6309 3836 6373 3840
rect 6309 3780 6313 3836
rect 6313 3780 6369 3836
rect 6369 3780 6373 3836
rect 6309 3776 6373 3780
rect 8116 3836 8180 3840
rect 8116 3780 8120 3836
rect 8120 3780 8176 3836
rect 8176 3780 8180 3836
rect 8116 3776 8180 3780
rect 8196 3836 8260 3840
rect 8196 3780 8200 3836
rect 8200 3780 8256 3836
rect 8256 3780 8260 3836
rect 8196 3776 8260 3780
rect 8276 3836 8340 3840
rect 8276 3780 8280 3836
rect 8280 3780 8336 3836
rect 8336 3780 8340 3836
rect 8276 3776 8340 3780
rect 8356 3836 8420 3840
rect 8356 3780 8360 3836
rect 8360 3780 8416 3836
rect 8416 3780 8420 3836
rect 8356 3776 8420 3780
rect 2635 3292 2699 3296
rect 2635 3236 2639 3292
rect 2639 3236 2695 3292
rect 2695 3236 2699 3292
rect 2635 3232 2699 3236
rect 2715 3292 2779 3296
rect 2715 3236 2719 3292
rect 2719 3236 2775 3292
rect 2775 3236 2779 3292
rect 2715 3232 2779 3236
rect 2795 3292 2859 3296
rect 2795 3236 2799 3292
rect 2799 3236 2855 3292
rect 2855 3236 2859 3292
rect 2795 3232 2859 3236
rect 2875 3292 2939 3296
rect 2875 3236 2879 3292
rect 2879 3236 2935 3292
rect 2935 3236 2939 3292
rect 2875 3232 2939 3236
rect 4682 3292 4746 3296
rect 4682 3236 4686 3292
rect 4686 3236 4742 3292
rect 4742 3236 4746 3292
rect 4682 3232 4746 3236
rect 4762 3292 4826 3296
rect 4762 3236 4766 3292
rect 4766 3236 4822 3292
rect 4822 3236 4826 3292
rect 4762 3232 4826 3236
rect 4842 3292 4906 3296
rect 4842 3236 4846 3292
rect 4846 3236 4902 3292
rect 4902 3236 4906 3292
rect 4842 3232 4906 3236
rect 4922 3292 4986 3296
rect 4922 3236 4926 3292
rect 4926 3236 4982 3292
rect 4982 3236 4986 3292
rect 4922 3232 4986 3236
rect 6729 3292 6793 3296
rect 6729 3236 6733 3292
rect 6733 3236 6789 3292
rect 6789 3236 6793 3292
rect 6729 3232 6793 3236
rect 6809 3292 6873 3296
rect 6809 3236 6813 3292
rect 6813 3236 6869 3292
rect 6869 3236 6873 3292
rect 6809 3232 6873 3236
rect 6889 3292 6953 3296
rect 6889 3236 6893 3292
rect 6893 3236 6949 3292
rect 6949 3236 6953 3292
rect 6889 3232 6953 3236
rect 6969 3292 7033 3296
rect 6969 3236 6973 3292
rect 6973 3236 7029 3292
rect 7029 3236 7033 3292
rect 6969 3232 7033 3236
rect 8776 3292 8840 3296
rect 8776 3236 8780 3292
rect 8780 3236 8836 3292
rect 8836 3236 8840 3292
rect 8776 3232 8840 3236
rect 8856 3292 8920 3296
rect 8856 3236 8860 3292
rect 8860 3236 8916 3292
rect 8916 3236 8920 3292
rect 8856 3232 8920 3236
rect 8936 3292 9000 3296
rect 8936 3236 8940 3292
rect 8940 3236 8996 3292
rect 8996 3236 9000 3292
rect 8936 3232 9000 3236
rect 9016 3292 9080 3296
rect 9016 3236 9020 3292
rect 9020 3236 9076 3292
rect 9076 3236 9080 3292
rect 9016 3232 9080 3236
rect 1975 2748 2039 2752
rect 1975 2692 1979 2748
rect 1979 2692 2035 2748
rect 2035 2692 2039 2748
rect 1975 2688 2039 2692
rect 2055 2748 2119 2752
rect 2055 2692 2059 2748
rect 2059 2692 2115 2748
rect 2115 2692 2119 2748
rect 2055 2688 2119 2692
rect 2135 2748 2199 2752
rect 2135 2692 2139 2748
rect 2139 2692 2195 2748
rect 2195 2692 2199 2748
rect 2135 2688 2199 2692
rect 2215 2748 2279 2752
rect 2215 2692 2219 2748
rect 2219 2692 2275 2748
rect 2275 2692 2279 2748
rect 2215 2688 2279 2692
rect 4022 2748 4086 2752
rect 4022 2692 4026 2748
rect 4026 2692 4082 2748
rect 4082 2692 4086 2748
rect 4022 2688 4086 2692
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 6069 2748 6133 2752
rect 6069 2692 6073 2748
rect 6073 2692 6129 2748
rect 6129 2692 6133 2748
rect 6069 2688 6133 2692
rect 6149 2748 6213 2752
rect 6149 2692 6153 2748
rect 6153 2692 6209 2748
rect 6209 2692 6213 2748
rect 6149 2688 6213 2692
rect 6229 2748 6293 2752
rect 6229 2692 6233 2748
rect 6233 2692 6289 2748
rect 6289 2692 6293 2748
rect 6229 2688 6293 2692
rect 6309 2748 6373 2752
rect 6309 2692 6313 2748
rect 6313 2692 6369 2748
rect 6369 2692 6373 2748
rect 6309 2688 6373 2692
rect 8116 2748 8180 2752
rect 8116 2692 8120 2748
rect 8120 2692 8176 2748
rect 8176 2692 8180 2748
rect 8116 2688 8180 2692
rect 8196 2748 8260 2752
rect 8196 2692 8200 2748
rect 8200 2692 8256 2748
rect 8256 2692 8260 2748
rect 8196 2688 8260 2692
rect 8276 2748 8340 2752
rect 8276 2692 8280 2748
rect 8280 2692 8336 2748
rect 8336 2692 8340 2748
rect 8276 2688 8340 2692
rect 8356 2748 8420 2752
rect 8356 2692 8360 2748
rect 8360 2692 8416 2748
rect 8416 2692 8420 2748
rect 8356 2688 8420 2692
rect 2635 2204 2699 2208
rect 2635 2148 2639 2204
rect 2639 2148 2695 2204
rect 2695 2148 2699 2204
rect 2635 2144 2699 2148
rect 2715 2204 2779 2208
rect 2715 2148 2719 2204
rect 2719 2148 2775 2204
rect 2775 2148 2779 2204
rect 2715 2144 2779 2148
rect 2795 2204 2859 2208
rect 2795 2148 2799 2204
rect 2799 2148 2855 2204
rect 2855 2148 2859 2204
rect 2795 2144 2859 2148
rect 2875 2204 2939 2208
rect 2875 2148 2879 2204
rect 2879 2148 2935 2204
rect 2935 2148 2939 2204
rect 2875 2144 2939 2148
rect 4682 2204 4746 2208
rect 4682 2148 4686 2204
rect 4686 2148 4742 2204
rect 4742 2148 4746 2204
rect 4682 2144 4746 2148
rect 4762 2204 4826 2208
rect 4762 2148 4766 2204
rect 4766 2148 4822 2204
rect 4822 2148 4826 2204
rect 4762 2144 4826 2148
rect 4842 2204 4906 2208
rect 4842 2148 4846 2204
rect 4846 2148 4902 2204
rect 4902 2148 4906 2204
rect 4842 2144 4906 2148
rect 4922 2204 4986 2208
rect 4922 2148 4926 2204
rect 4926 2148 4982 2204
rect 4982 2148 4986 2204
rect 4922 2144 4986 2148
rect 6729 2204 6793 2208
rect 6729 2148 6733 2204
rect 6733 2148 6789 2204
rect 6789 2148 6793 2204
rect 6729 2144 6793 2148
rect 6809 2204 6873 2208
rect 6809 2148 6813 2204
rect 6813 2148 6869 2204
rect 6869 2148 6873 2204
rect 6809 2144 6873 2148
rect 6889 2204 6953 2208
rect 6889 2148 6893 2204
rect 6893 2148 6949 2204
rect 6949 2148 6953 2204
rect 6889 2144 6953 2148
rect 6969 2204 7033 2208
rect 6969 2148 6973 2204
rect 6973 2148 7029 2204
rect 7029 2148 7033 2204
rect 6969 2144 7033 2148
rect 8776 2204 8840 2208
rect 8776 2148 8780 2204
rect 8780 2148 8836 2204
rect 8836 2148 8840 2204
rect 8776 2144 8840 2148
rect 8856 2204 8920 2208
rect 8856 2148 8860 2204
rect 8860 2148 8916 2204
rect 8916 2148 8920 2204
rect 8856 2144 8920 2148
rect 8936 2204 9000 2208
rect 8936 2148 8940 2204
rect 8940 2148 8996 2204
rect 8996 2148 9000 2204
rect 8936 2144 9000 2148
rect 9016 2204 9080 2208
rect 9016 2148 9020 2204
rect 9020 2148 9076 2204
rect 9076 2148 9080 2204
rect 9016 2144 9080 2148
<< metal4 >>
rect 1967 10368 2287 10384
rect 1967 10304 1975 10368
rect 2039 10304 2055 10368
rect 2119 10304 2135 10368
rect 2199 10304 2215 10368
rect 2279 10304 2287 10368
rect 1967 9434 2287 10304
rect 1967 9280 2009 9434
rect 2245 9280 2287 9434
rect 1967 9216 1975 9280
rect 2279 9216 2287 9280
rect 1967 9198 2009 9216
rect 2245 9198 2287 9216
rect 1967 8192 2287 9198
rect 1967 8128 1975 8192
rect 2039 8128 2055 8192
rect 2119 8128 2135 8192
rect 2199 8128 2215 8192
rect 2279 8128 2287 8192
rect 1967 7394 2287 8128
rect 1967 7158 2009 7394
rect 2245 7158 2287 7394
rect 1967 7104 2287 7158
rect 1967 7040 1975 7104
rect 2039 7040 2055 7104
rect 2119 7040 2135 7104
rect 2199 7040 2215 7104
rect 2279 7040 2287 7104
rect 1967 6016 2287 7040
rect 1967 5952 1975 6016
rect 2039 5952 2055 6016
rect 2119 5952 2135 6016
rect 2199 5952 2215 6016
rect 2279 5952 2287 6016
rect 1967 5354 2287 5952
rect 1967 5118 2009 5354
rect 2245 5118 2287 5354
rect 1967 4928 2287 5118
rect 1967 4864 1975 4928
rect 2039 4864 2055 4928
rect 2119 4864 2135 4928
rect 2199 4864 2215 4928
rect 2279 4864 2287 4928
rect 1967 3840 2287 4864
rect 1967 3776 1975 3840
rect 2039 3776 2055 3840
rect 2119 3776 2135 3840
rect 2199 3776 2215 3840
rect 2279 3776 2287 3840
rect 1967 3314 2287 3776
rect 1967 3078 2009 3314
rect 2245 3078 2287 3314
rect 1967 2752 2287 3078
rect 1967 2688 1975 2752
rect 2039 2688 2055 2752
rect 2119 2688 2135 2752
rect 2199 2688 2215 2752
rect 2279 2688 2287 2752
rect 1967 2128 2287 2688
rect 2627 10094 2947 10384
rect 2627 9858 2669 10094
rect 2905 9858 2947 10094
rect 2627 9824 2947 9858
rect 2627 9760 2635 9824
rect 2699 9760 2715 9824
rect 2779 9760 2795 9824
rect 2859 9760 2875 9824
rect 2939 9760 2947 9824
rect 2627 8736 2947 9760
rect 2627 8672 2635 8736
rect 2699 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2875 8736
rect 2939 8672 2947 8736
rect 2627 8054 2947 8672
rect 2627 7818 2669 8054
rect 2905 7818 2947 8054
rect 2627 7648 2947 7818
rect 2627 7584 2635 7648
rect 2699 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2875 7648
rect 2939 7584 2947 7648
rect 2627 6560 2947 7584
rect 2627 6496 2635 6560
rect 2699 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2875 6560
rect 2939 6496 2947 6560
rect 2627 6014 2947 6496
rect 2627 5778 2669 6014
rect 2905 5778 2947 6014
rect 2627 5472 2947 5778
rect 2627 5408 2635 5472
rect 2699 5408 2715 5472
rect 2779 5408 2795 5472
rect 2859 5408 2875 5472
rect 2939 5408 2947 5472
rect 2627 4384 2947 5408
rect 2627 4320 2635 4384
rect 2699 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2875 4384
rect 2939 4320 2947 4384
rect 2627 3974 2947 4320
rect 2627 3738 2669 3974
rect 2905 3738 2947 3974
rect 2627 3296 2947 3738
rect 2627 3232 2635 3296
rect 2699 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2875 3296
rect 2939 3232 2947 3296
rect 2627 2208 2947 3232
rect 2627 2144 2635 2208
rect 2699 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2875 2208
rect 2939 2144 2947 2208
rect 2627 2128 2947 2144
rect 4014 10368 4334 10384
rect 4014 10304 4022 10368
rect 4086 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4334 10368
rect 4014 9434 4334 10304
rect 4014 9280 4056 9434
rect 4292 9280 4334 9434
rect 4014 9216 4022 9280
rect 4326 9216 4334 9280
rect 4014 9198 4056 9216
rect 4292 9198 4334 9216
rect 4014 8192 4334 9198
rect 4014 8128 4022 8192
rect 4086 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4334 8192
rect 4014 7394 4334 8128
rect 4014 7158 4056 7394
rect 4292 7158 4334 7394
rect 4014 7104 4334 7158
rect 4014 7040 4022 7104
rect 4086 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4334 7104
rect 4014 6016 4334 7040
rect 4014 5952 4022 6016
rect 4086 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4334 6016
rect 4014 5354 4334 5952
rect 4014 5118 4056 5354
rect 4292 5118 4334 5354
rect 4014 4928 4334 5118
rect 4014 4864 4022 4928
rect 4086 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4334 4928
rect 4014 3840 4334 4864
rect 4014 3776 4022 3840
rect 4086 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4334 3840
rect 4014 3314 4334 3776
rect 4014 3078 4056 3314
rect 4292 3078 4334 3314
rect 4014 2752 4334 3078
rect 4014 2688 4022 2752
rect 4086 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4334 2752
rect 4014 2128 4334 2688
rect 4674 10094 4994 10384
rect 4674 9858 4716 10094
rect 4952 9858 4994 10094
rect 4674 9824 4994 9858
rect 4674 9760 4682 9824
rect 4746 9760 4762 9824
rect 4826 9760 4842 9824
rect 4906 9760 4922 9824
rect 4986 9760 4994 9824
rect 4674 8736 4994 9760
rect 4674 8672 4682 8736
rect 4746 8672 4762 8736
rect 4826 8672 4842 8736
rect 4906 8672 4922 8736
rect 4986 8672 4994 8736
rect 4674 8054 4994 8672
rect 4674 7818 4716 8054
rect 4952 7818 4994 8054
rect 4674 7648 4994 7818
rect 4674 7584 4682 7648
rect 4746 7584 4762 7648
rect 4826 7584 4842 7648
rect 4906 7584 4922 7648
rect 4986 7584 4994 7648
rect 4674 6560 4994 7584
rect 4674 6496 4682 6560
rect 4746 6496 4762 6560
rect 4826 6496 4842 6560
rect 4906 6496 4922 6560
rect 4986 6496 4994 6560
rect 4674 6014 4994 6496
rect 4674 5778 4716 6014
rect 4952 5778 4994 6014
rect 4674 5472 4994 5778
rect 4674 5408 4682 5472
rect 4746 5408 4762 5472
rect 4826 5408 4842 5472
rect 4906 5408 4922 5472
rect 4986 5408 4994 5472
rect 4674 4384 4994 5408
rect 4674 4320 4682 4384
rect 4746 4320 4762 4384
rect 4826 4320 4842 4384
rect 4906 4320 4922 4384
rect 4986 4320 4994 4384
rect 4674 3974 4994 4320
rect 4674 3738 4716 3974
rect 4952 3738 4994 3974
rect 4674 3296 4994 3738
rect 4674 3232 4682 3296
rect 4746 3232 4762 3296
rect 4826 3232 4842 3296
rect 4906 3232 4922 3296
rect 4986 3232 4994 3296
rect 4674 2208 4994 3232
rect 4674 2144 4682 2208
rect 4746 2144 4762 2208
rect 4826 2144 4842 2208
rect 4906 2144 4922 2208
rect 4986 2144 4994 2208
rect 4674 2128 4994 2144
rect 6061 10368 6381 10384
rect 6061 10304 6069 10368
rect 6133 10304 6149 10368
rect 6213 10304 6229 10368
rect 6293 10304 6309 10368
rect 6373 10304 6381 10368
rect 6061 9434 6381 10304
rect 6061 9280 6103 9434
rect 6339 9280 6381 9434
rect 6061 9216 6069 9280
rect 6373 9216 6381 9280
rect 6061 9198 6103 9216
rect 6339 9198 6381 9216
rect 6061 8192 6381 9198
rect 6061 8128 6069 8192
rect 6133 8128 6149 8192
rect 6213 8128 6229 8192
rect 6293 8128 6309 8192
rect 6373 8128 6381 8192
rect 6061 7394 6381 8128
rect 6061 7158 6103 7394
rect 6339 7158 6381 7394
rect 6061 7104 6381 7158
rect 6061 7040 6069 7104
rect 6133 7040 6149 7104
rect 6213 7040 6229 7104
rect 6293 7040 6309 7104
rect 6373 7040 6381 7104
rect 6061 6016 6381 7040
rect 6061 5952 6069 6016
rect 6133 5952 6149 6016
rect 6213 5952 6229 6016
rect 6293 5952 6309 6016
rect 6373 5952 6381 6016
rect 6061 5354 6381 5952
rect 6061 5118 6103 5354
rect 6339 5118 6381 5354
rect 6061 4928 6381 5118
rect 6061 4864 6069 4928
rect 6133 4864 6149 4928
rect 6213 4864 6229 4928
rect 6293 4864 6309 4928
rect 6373 4864 6381 4928
rect 6061 3840 6381 4864
rect 6061 3776 6069 3840
rect 6133 3776 6149 3840
rect 6213 3776 6229 3840
rect 6293 3776 6309 3840
rect 6373 3776 6381 3840
rect 6061 3314 6381 3776
rect 6061 3078 6103 3314
rect 6339 3078 6381 3314
rect 6061 2752 6381 3078
rect 6061 2688 6069 2752
rect 6133 2688 6149 2752
rect 6213 2688 6229 2752
rect 6293 2688 6309 2752
rect 6373 2688 6381 2752
rect 6061 2128 6381 2688
rect 6721 10094 7041 10384
rect 6721 9858 6763 10094
rect 6999 9858 7041 10094
rect 6721 9824 7041 9858
rect 6721 9760 6729 9824
rect 6793 9760 6809 9824
rect 6873 9760 6889 9824
rect 6953 9760 6969 9824
rect 7033 9760 7041 9824
rect 6721 8736 7041 9760
rect 6721 8672 6729 8736
rect 6793 8672 6809 8736
rect 6873 8672 6889 8736
rect 6953 8672 6969 8736
rect 7033 8672 7041 8736
rect 6721 8054 7041 8672
rect 6721 7818 6763 8054
rect 6999 7818 7041 8054
rect 6721 7648 7041 7818
rect 6721 7584 6729 7648
rect 6793 7584 6809 7648
rect 6873 7584 6889 7648
rect 6953 7584 6969 7648
rect 7033 7584 7041 7648
rect 6721 6560 7041 7584
rect 6721 6496 6729 6560
rect 6793 6496 6809 6560
rect 6873 6496 6889 6560
rect 6953 6496 6969 6560
rect 7033 6496 7041 6560
rect 6721 6014 7041 6496
rect 6721 5778 6763 6014
rect 6999 5778 7041 6014
rect 6721 5472 7041 5778
rect 6721 5408 6729 5472
rect 6793 5408 6809 5472
rect 6873 5408 6889 5472
rect 6953 5408 6969 5472
rect 7033 5408 7041 5472
rect 6721 4384 7041 5408
rect 6721 4320 6729 4384
rect 6793 4320 6809 4384
rect 6873 4320 6889 4384
rect 6953 4320 6969 4384
rect 7033 4320 7041 4384
rect 6721 3974 7041 4320
rect 6721 3738 6763 3974
rect 6999 3738 7041 3974
rect 6721 3296 7041 3738
rect 6721 3232 6729 3296
rect 6793 3232 6809 3296
rect 6873 3232 6889 3296
rect 6953 3232 6969 3296
rect 7033 3232 7041 3296
rect 6721 2208 7041 3232
rect 6721 2144 6729 2208
rect 6793 2144 6809 2208
rect 6873 2144 6889 2208
rect 6953 2144 6969 2208
rect 7033 2144 7041 2208
rect 6721 2128 7041 2144
rect 8108 10368 8428 10384
rect 8108 10304 8116 10368
rect 8180 10304 8196 10368
rect 8260 10304 8276 10368
rect 8340 10304 8356 10368
rect 8420 10304 8428 10368
rect 8108 9434 8428 10304
rect 8108 9280 8150 9434
rect 8386 9280 8428 9434
rect 8108 9216 8116 9280
rect 8420 9216 8428 9280
rect 8108 9198 8150 9216
rect 8386 9198 8428 9216
rect 8108 8192 8428 9198
rect 8108 8128 8116 8192
rect 8180 8128 8196 8192
rect 8260 8128 8276 8192
rect 8340 8128 8356 8192
rect 8420 8128 8428 8192
rect 8108 7394 8428 8128
rect 8108 7158 8150 7394
rect 8386 7158 8428 7394
rect 8108 7104 8428 7158
rect 8108 7040 8116 7104
rect 8180 7040 8196 7104
rect 8260 7040 8276 7104
rect 8340 7040 8356 7104
rect 8420 7040 8428 7104
rect 8108 6016 8428 7040
rect 8108 5952 8116 6016
rect 8180 5952 8196 6016
rect 8260 5952 8276 6016
rect 8340 5952 8356 6016
rect 8420 5952 8428 6016
rect 8108 5354 8428 5952
rect 8108 5118 8150 5354
rect 8386 5118 8428 5354
rect 8108 4928 8428 5118
rect 8108 4864 8116 4928
rect 8180 4864 8196 4928
rect 8260 4864 8276 4928
rect 8340 4864 8356 4928
rect 8420 4864 8428 4928
rect 8108 3840 8428 4864
rect 8108 3776 8116 3840
rect 8180 3776 8196 3840
rect 8260 3776 8276 3840
rect 8340 3776 8356 3840
rect 8420 3776 8428 3840
rect 8108 3314 8428 3776
rect 8108 3078 8150 3314
rect 8386 3078 8428 3314
rect 8108 2752 8428 3078
rect 8108 2688 8116 2752
rect 8180 2688 8196 2752
rect 8260 2688 8276 2752
rect 8340 2688 8356 2752
rect 8420 2688 8428 2752
rect 8108 2128 8428 2688
rect 8768 10094 9088 10384
rect 8768 9858 8810 10094
rect 9046 9858 9088 10094
rect 8768 9824 9088 9858
rect 8768 9760 8776 9824
rect 8840 9760 8856 9824
rect 8920 9760 8936 9824
rect 9000 9760 9016 9824
rect 9080 9760 9088 9824
rect 8768 8736 9088 9760
rect 8768 8672 8776 8736
rect 8840 8672 8856 8736
rect 8920 8672 8936 8736
rect 9000 8672 9016 8736
rect 9080 8672 9088 8736
rect 8768 8054 9088 8672
rect 8768 7818 8810 8054
rect 9046 7818 9088 8054
rect 8768 7648 9088 7818
rect 8768 7584 8776 7648
rect 8840 7584 8856 7648
rect 8920 7584 8936 7648
rect 9000 7584 9016 7648
rect 9080 7584 9088 7648
rect 8768 6560 9088 7584
rect 8768 6496 8776 6560
rect 8840 6496 8856 6560
rect 8920 6496 8936 6560
rect 9000 6496 9016 6560
rect 9080 6496 9088 6560
rect 8768 6014 9088 6496
rect 8768 5778 8810 6014
rect 9046 5778 9088 6014
rect 8768 5472 9088 5778
rect 8768 5408 8776 5472
rect 8840 5408 8856 5472
rect 8920 5408 8936 5472
rect 9000 5408 9016 5472
rect 9080 5408 9088 5472
rect 8768 4384 9088 5408
rect 8768 4320 8776 4384
rect 8840 4320 8856 4384
rect 8920 4320 8936 4384
rect 9000 4320 9016 4384
rect 9080 4320 9088 4384
rect 8768 3974 9088 4320
rect 8768 3738 8810 3974
rect 9046 3738 9088 3974
rect 8768 3296 9088 3738
rect 8768 3232 8776 3296
rect 8840 3232 8856 3296
rect 8920 3232 8936 3296
rect 9000 3232 9016 3296
rect 9080 3232 9088 3296
rect 8768 2208 9088 3232
rect 8768 2144 8776 2208
rect 8840 2144 8856 2208
rect 8920 2144 8936 2208
rect 9000 2144 9016 2208
rect 9080 2144 9088 2208
rect 8768 2128 9088 2144
<< via4 >>
rect 2009 9280 2245 9434
rect 2009 9216 2039 9280
rect 2039 9216 2055 9280
rect 2055 9216 2119 9280
rect 2119 9216 2135 9280
rect 2135 9216 2199 9280
rect 2199 9216 2215 9280
rect 2215 9216 2245 9280
rect 2009 9198 2245 9216
rect 2009 7158 2245 7394
rect 2009 5118 2245 5354
rect 2009 3078 2245 3314
rect 2669 9858 2905 10094
rect 2669 7818 2905 8054
rect 2669 5778 2905 6014
rect 2669 3738 2905 3974
rect 4056 9280 4292 9434
rect 4056 9216 4086 9280
rect 4086 9216 4102 9280
rect 4102 9216 4166 9280
rect 4166 9216 4182 9280
rect 4182 9216 4246 9280
rect 4246 9216 4262 9280
rect 4262 9216 4292 9280
rect 4056 9198 4292 9216
rect 4056 7158 4292 7394
rect 4056 5118 4292 5354
rect 4056 3078 4292 3314
rect 4716 9858 4952 10094
rect 4716 7818 4952 8054
rect 4716 5778 4952 6014
rect 4716 3738 4952 3974
rect 6103 9280 6339 9434
rect 6103 9216 6133 9280
rect 6133 9216 6149 9280
rect 6149 9216 6213 9280
rect 6213 9216 6229 9280
rect 6229 9216 6293 9280
rect 6293 9216 6309 9280
rect 6309 9216 6339 9280
rect 6103 9198 6339 9216
rect 6103 7158 6339 7394
rect 6103 5118 6339 5354
rect 6103 3078 6339 3314
rect 6763 9858 6999 10094
rect 6763 7818 6999 8054
rect 6763 5778 6999 6014
rect 6763 3738 6999 3974
rect 8150 9280 8386 9434
rect 8150 9216 8180 9280
rect 8180 9216 8196 9280
rect 8196 9216 8260 9280
rect 8260 9216 8276 9280
rect 8276 9216 8340 9280
rect 8340 9216 8356 9280
rect 8356 9216 8386 9280
rect 8150 9198 8386 9216
rect 8150 7158 8386 7394
rect 8150 5118 8386 5354
rect 8150 3078 8386 3314
rect 8810 9858 9046 10094
rect 8810 7818 9046 8054
rect 8810 5778 9046 6014
rect 8810 3738 9046 3974
<< metal5 >>
rect 1056 10094 9340 10136
rect 1056 9858 2669 10094
rect 2905 9858 4716 10094
rect 4952 9858 6763 10094
rect 6999 9858 8810 10094
rect 9046 9858 9340 10094
rect 1056 9816 9340 9858
rect 1056 9434 9340 9476
rect 1056 9198 2009 9434
rect 2245 9198 4056 9434
rect 4292 9198 6103 9434
rect 6339 9198 8150 9434
rect 8386 9198 9340 9434
rect 1056 9156 9340 9198
rect 1056 8054 9340 8096
rect 1056 7818 2669 8054
rect 2905 7818 4716 8054
rect 4952 7818 6763 8054
rect 6999 7818 8810 8054
rect 9046 7818 9340 8054
rect 1056 7776 9340 7818
rect 1056 7394 9340 7436
rect 1056 7158 2009 7394
rect 2245 7158 4056 7394
rect 4292 7158 6103 7394
rect 6339 7158 8150 7394
rect 8386 7158 9340 7394
rect 1056 7116 9340 7158
rect 1056 6014 9340 6056
rect 1056 5778 2669 6014
rect 2905 5778 4716 6014
rect 4952 5778 6763 6014
rect 6999 5778 8810 6014
rect 9046 5778 9340 6014
rect 1056 5736 9340 5778
rect 1056 5354 9340 5396
rect 1056 5118 2009 5354
rect 2245 5118 4056 5354
rect 4292 5118 6103 5354
rect 6339 5118 8150 5354
rect 8386 5118 9340 5354
rect 1056 5076 9340 5118
rect 1056 3974 9340 4016
rect 1056 3738 2669 3974
rect 2905 3738 4716 3974
rect 4952 3738 6763 3974
rect 6999 3738 8810 3974
rect 9046 3738 9340 3974
rect 1056 3696 9340 3738
rect 1056 3314 9340 3356
rect 1056 3078 2009 3314
rect 2245 3078 4056 3314
rect 4292 3078 6103 3314
rect 6339 3078 8150 3314
rect 8386 3078 9340 3314
rect 1056 3036 9340 3078
use sky130_fd_sc_hd__buf_2  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1723858470
transform -1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_2  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5336 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6256 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1840 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2576 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4968 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2392 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _074_
timestamp 1723858470
transform 1 0 5520 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _076_
timestamp 1723858470
transform 1 0 5520 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_1  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7084 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7544 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _083_
timestamp 1723858470
transform 1 0 7636 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _084_
timestamp 1723858470
transform -1 0 8740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _085_
timestamp 1723858470
transform -1 0 8648 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _086_
timestamp 1723858470
transform -1 0 8740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8188 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _089_
timestamp 1723858470
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3404 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _091_
timestamp 1723858470
transform 1 0 3404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _092_
timestamp 1723858470
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand4b_1  _094_
timestamp 1723858470
transform 1 0 1932 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6808 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7360 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _097_
timestamp 1723858470
transform -1 0 8372 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _098_
timestamp 1723858470
transform -1 0 8832 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _102_
timestamp 1723858470
transform 1 0 2576 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _103_
timestamp 1723858470
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _104_
timestamp 1723858470
transform -1 0 4416 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _105_
timestamp 1723858470
transform -1 0 4416 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _106_
timestamp 1723858470
transform -1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _107_
timestamp 1723858470
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _108_
timestamp 1723858470
transform 1 0 2944 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _110_
timestamp 1723858470
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _111_
timestamp 1723858470
transform -1 0 6992 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _112_
timestamp 1723858470
transform 1 0 6992 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _113_
timestamp 1723858470
transform -1 0 6808 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _115_
timestamp 1723858470
transform 1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5428 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5336 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3956 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _120_
timestamp 1723858470
transform 1 0 5244 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _122_
timestamp 1723858470
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _123_
timestamp 1723858470
transform 1 0 5152 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7176 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _125_
timestamp 1723858470
transform -1 0 2852 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _126_
timestamp 1723858470
transform -1 0 2852 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _127_
timestamp 1723858470
transform 1 0 7544 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1723858470
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1723858470
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_36
timestamp 1723858470
transform 1 0 4416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_44
timestamp 1723858470
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48
timestamp 1723858470
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_76
timestamp 1723858470
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1723858470
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_7
timestamp 1723858470
transform 1 0 1748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 1723858470
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_40
timestamp 1723858470
transform 1 0 4784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1723858470
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_9
timestamp 1723858470
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_13
timestamp 1723858470
transform 1 0 2300 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_46
timestamp 1723858470
transform 1 0 5336 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_55
timestamp 1723858470
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_67
timestamp 1723858470
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_79
timestamp 1723858470
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1723858470
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1723858470
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1723858470
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1723858470
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_39
timestamp 1723858470
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_47
timestamp 1723858470
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_64
timestamp 1723858470
transform 1 0 6992 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_76
timestamp 1723858470
transform 1 0 8096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_84
timestamp 1723858470
transform 1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1723858470
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1723858470
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1723858470
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_40
timestamp 1723858470
transform 1 0 4784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_48
timestamp 1723858470
transform 1 0 5520 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_56
timestamp 1723858470
transform 1 0 6256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_68
timestamp 1723858470
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 1723858470
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1723858470
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1723858470
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_7
timestamp 1723858470
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_15
timestamp 1723858470
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_29
timestamp 1723858470
transform 1 0 3772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_41
timestamp 1723858470
transform 1 0 4876 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1723858470
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_69
timestamp 1723858470
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_83
timestamp 1723858470
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_9
timestamp 1723858470
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1723858470
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_40
timestamp 1723858470
transform 1 0 4784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_74
timestamp 1723858470
transform 1 0 7912 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_80
timestamp 1723858470
transform 1 0 8464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1723858470
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 1723858470
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_21
timestamp 1723858470
transform 1 0 3036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_27
timestamp 1723858470
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_36
timestamp 1723858470
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1723858470
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1723858470
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1723858470
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_69
timestamp 1723858470
transform 1 0 7452 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_82
timestamp 1723858470
transform 1 0 8648 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1723858470
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_15
timestamp 1723858470
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_19
timestamp 1723858470
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_24
timestamp 1723858470
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_39
timestamp 1723858470
transform 1 0 4692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_47
timestamp 1723858470
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_52
timestamp 1723858470
transform 1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_60
timestamp 1723858470
transform 1 0 6624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1723858470
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 1723858470
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_36
timestamp 1723858470
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_44
timestamp 1723858470
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1723858470
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_64
timestamp 1723858470
transform 1 0 6992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_70
timestamp 1723858470
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_76
timestamp 1723858470
transform 1 0 8096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_84
timestamp 1723858470
transform 1 0 8832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_19
timestamp 1723858470
transform 1 0 2852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1723858470
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_33
timestamp 1723858470
transform 1 0 4140 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 1723858470
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_51
timestamp 1723858470
transform 1 0 5796 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_63
timestamp 1723858470
transform 1 0 6900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_75
timestamp 1723858470
transform 1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_79
timestamp 1723858470
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1723858470
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_7
timestamp 1723858470
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_19
timestamp 1723858470
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_31
timestamp 1723858470
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_43
timestamp 1723858470
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1723858470
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1723858470
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1723858470
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1723858470
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_15
timestamp 1723858470
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_23
timestamp 1723858470
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1723858470
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1723858470
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_37
timestamp 1723858470
transform 1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_55
timestamp 1723858470
transform 1 0 6164 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_67
timestamp 1723858470
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_73
timestamp 1723858470
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1723858470
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1723858470
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1723858470
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_15
timestamp 1723858470
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_30
timestamp 1723858470
transform 1 0 3864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_36
timestamp 1723858470
transform 1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_42
timestamp 1723858470
transform 1 0 4968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_48
timestamp 1723858470
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_52
timestamp 1723858470
transform 1 0 5888 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_62
timestamp 1723858470
transform 1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_70
timestamp 1723858470
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_84
timestamp 1723858470
transform 1 0 8832 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_10
timestamp 1723858470
transform 1 0 2024 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_22
timestamp 1723858470
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_35
timestamp 1723858470
transform 1 0 4324 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_47
timestamp 1723858470
transform 1 0 5428 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_55
timestamp 1723858470
transform 1 0 6164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_57
timestamp 1723858470
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_63
timestamp 1723858470
transform 1 0 6900 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_71
timestamp 1723858470
transform 1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1723858470
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1723858470
transform -1 0 8832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1723858470
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1723858470
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1723858470
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1723858470
transform 1 0 3956 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1723858470
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1723858470
transform -1 0 8832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1723858470
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1723858470
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1723858470
transform 1 0 1748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1723858470
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1723858470
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1723858470
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1723858470
transform -1 0 8464 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1723858470
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1723858470
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1723858470
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1723858470
transform -1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1723858470
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1723858470
transform -1 0 9292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1723858470
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1723858470
transform -1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1723858470
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1723858470
transform -1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1723858470
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1723858470
transform -1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1723858470
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1723858470
transform -1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1723858470
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1723858470
transform -1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1723858470
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1723858470
transform -1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1723858470
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1723858470
transform -1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1723858470
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1723858470
transform -1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1723858470
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1723858470
transform -1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1723858470
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1723858470
transform -1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1723858470
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1723858470
transform -1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1723858470
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1723858470
transform -1 0 9292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1723858470
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1723858470
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1723858470
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1723858470
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1723858470
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1723858470
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1723858470
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1723858470
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1723858470
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1723858470
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1723858470
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1723858470
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1723858470
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1723858470
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1723858470
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1723858470
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1723858470
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1723858470
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1723858470
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1723858470
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1723858470
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1723858470
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1723858470
transform 1 0 6256 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1723858470
transform 1 0 8832 0 1 9792
box -38 -48 130 592
<< labels >>
flabel metal3 s 9673 8168 10473 8288 0 FreeSans 480 0 0 0 A[0]
port 0 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 A[1]
port 1 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 A[2]
port 2 nsew signal input
flabel metal2 s 6458 11817 6514 12617 0 FreeSans 224 90 0 0 A[3]
port 3 nsew signal input
flabel metal2 s 3882 11817 3938 12617 0 FreeSans 224 90 0 0 B[0]
port 4 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 B[1]
port 5 nsew signal input
flabel metal3 s 9673 10888 10473 11008 0 FreeSans 480 0 0 0 B[2]
port 6 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 B[3]
port 7 nsew signal input
flabel metal4 s 2627 2128 2947 10384 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 4674 2128 4994 10384 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 6721 2128 7041 10384 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 8768 2128 9088 10384 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 3696 9340 4016 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 5736 9340 6056 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 7776 9340 8096 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 9816 9340 10136 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 1967 2128 2287 10384 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 4014 2128 4334 10384 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 6061 2128 6381 10384 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 8108 2128 8428 10384 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 3036 9340 3356 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 5076 9340 5396 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 7116 9340 7436 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 9156 9340 9476 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 clk
port 10 nsew signal input
flabel metal3 s 9673 2728 10473 2848 0 FreeSans 480 0 0 0 result[0]
port 11 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 result[1]
port 12 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 result[2]
port 13 nsew signal tristate
flabel metal2 s 9034 11817 9090 12617 0 FreeSans 224 90 0 0 result[3]
port 14 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 rst
port 15 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 sel[0]
port 16 nsew signal input
flabel metal2 s 1306 11817 1362 12617 0 FreeSans 224 90 0 0 sel[1]
port 17 nsew signal input
flabel metal3 s 9673 5448 10473 5568 0 FreeSans 480 0 0 0 sel[2]
port 18 nsew signal input
rlabel metal1 5198 9792 5198 9792 0 VGND
rlabel metal1 5198 10336 5198 10336 0 VPWR
rlabel metal1 8970 7854 8970 7854 0 A[0]
rlabel metal2 10350 1588 10350 1588 0 A[1]
rlabel metal3 820 10948 820 10948 0 A[2]
rlabel metal1 6578 10030 6578 10030 0 A[3]
rlabel metal1 4002 10030 4002 10030 0 B[0]
rlabel metal1 782 3026 782 3026 0 B[1]
rlabel metal1 8970 10030 8970 10030 0 B[2]
rlabel metal2 7774 1588 7774 1588 0 B[3]
rlabel metal1 7298 3094 7298 3094 0 _000_
rlabel metal1 3419 2346 3419 2346 0 _001_
rlabel metal1 3358 7888 3358 7888 0 _002_
rlabel metal1 6302 8058 6302 8058 0 _003_
rlabel metal1 4416 6698 4416 6698 0 _004_
rlabel metal1 4324 6766 4324 6766 0 _005_
rlabel metal2 5198 3672 5198 3672 0 _006_
rlabel metal1 6348 4794 6348 4794 0 _007_
rlabel metal2 4462 5134 4462 5134 0 _008_
rlabel metal1 6302 4046 6302 4046 0 _009_
rlabel metal1 5888 3570 5888 3570 0 _010_
rlabel metal1 2893 5168 2893 5168 0 _011_
rlabel metal1 4738 6222 4738 6222 0 _012_
rlabel metal1 5612 3706 5612 3706 0 _013_
rlabel metal1 2990 3434 2990 3434 0 _014_
rlabel metal1 3772 2278 3772 2278 0 _015_
rlabel metal2 5934 3094 5934 3094 0 _016_
rlabel metal1 6164 3094 6164 3094 0 _017_
rlabel metal1 6992 3010 6992 3010 0 _018_
rlabel metal2 3910 2587 3910 2587 0 _019_
rlabel metal1 3358 6630 3358 6630 0 _020_
rlabel metal1 7958 6800 7958 6800 0 _021_
rlabel metal1 8004 6970 8004 6970 0 _022_
rlabel metal1 8142 6766 8142 6766 0 _023_
rlabel metal1 8004 7174 8004 7174 0 _024_
rlabel metal1 8280 6290 8280 6290 0 _025_
rlabel metal2 7958 5678 7958 5678 0 _026_
rlabel metal1 7774 5134 7774 5134 0 _027_
rlabel metal1 4324 5202 4324 5202 0 _028_
rlabel metal1 4094 4658 4094 4658 0 _029_
rlabel metal1 3588 4794 3588 4794 0 _030_
rlabel metal1 2714 5304 2714 5304 0 _031_
rlabel metal1 3634 2414 3634 2414 0 _032_
rlabel metal1 4324 2618 4324 2618 0 _033_
rlabel metal2 2990 7616 2990 7616 0 _034_
rlabel metal1 5152 8942 5152 8942 0 _035_
rlabel metal1 8326 9588 8326 9588 0 _036_
rlabel metal1 4094 9588 4094 9588 0 _037_
rlabel metal1 4646 9350 4646 9350 0 _038_
rlabel metal1 2714 9588 2714 9588 0 _039_
rlabel metal1 4876 9554 4876 9554 0 _040_
rlabel metal1 2898 9078 2898 9078 0 _041_
rlabel metal1 2990 6800 2990 6800 0 _042_
rlabel metal1 4094 5712 4094 5712 0 _043_
rlabel metal1 4462 5882 4462 5882 0 _044_
rlabel metal1 3496 6426 3496 6426 0 _045_
rlabel metal1 3128 7854 3128 7854 0 _046_
rlabel metal1 3588 8058 3588 8058 0 _047_
rlabel metal1 4922 9452 4922 9452 0 _048_
rlabel metal1 5842 9010 5842 9010 0 _049_
rlabel metal1 5980 7514 5980 7514 0 _050_
rlabel metal1 6762 9520 6762 9520 0 _051_
rlabel metal1 5888 9554 5888 9554 0 _052_
rlabel metal1 5658 9588 5658 9588 0 _053_
rlabel metal1 4922 8976 4922 8976 0 _054_
rlabel metal1 6026 8874 6026 8874 0 _055_
rlabel metal1 5428 7718 5428 7718 0 _056_
rlabel metal1 5336 7514 5336 7514 0 _057_
rlabel metal1 5060 6290 5060 6290 0 _058_
rlabel metal1 5198 6222 5198 6222 0 _059_
rlabel metal2 5198 7106 5198 7106 0 _060_
rlabel metal2 5566 7514 5566 7514 0 _061_
rlabel metal2 2622 1367 2622 1367 0 clk
rlabel metal2 4370 5236 4370 5236 0 clknet_0_clk
rlabel metal1 3082 2924 3082 2924 0 clknet_1_0__leaf_clk
rlabel metal1 2806 7956 2806 7956 0 clknet_1_1__leaf_clk
rlabel metal2 8510 6392 8510 6392 0 net1
rlabel metal1 2162 7412 2162 7412 0 net10
rlabel metal1 1932 6290 1932 6290 0 net11
rlabel metal1 7222 5610 7222 5610 0 net12
rlabel metal1 8648 3026 8648 3026 0 net13
rlabel metal1 1472 2618 1472 2618 0 net14
rlabel metal1 1472 5678 1472 5678 0 net15
rlabel metal1 8740 8602 8740 8602 0 net16
rlabel metal1 8602 6766 8602 6766 0 net2
rlabel metal1 3266 9690 3266 9690 0 net3
rlabel metal1 6762 7412 6762 7412 0 net4
rlabel metal1 5704 9962 5704 9962 0 net5
rlabel metal2 7452 6834 7452 6834 0 net6
rlabel metal1 4738 5644 4738 5644 0 net7
rlabel metal2 7866 2689 7866 2689 0 net8
rlabel metal1 5566 2618 5566 2618 0 net9
rlabel via2 8878 2805 8878 2805 0 result[0]
rlabel metal3 820 2788 820 2788 0 result[1]
rlabel metal3 1142 5508 1142 5508 0 result[2]
rlabel metal1 8648 10234 8648 10234 0 result[3]
rlabel metal2 5198 1027 5198 1027 0 rst
rlabel metal3 1050 8228 1050 8228 0 sel[0]
rlabel metal1 1794 10064 1794 10064 0 sel[1]
rlabel metal1 9062 5678 9062 5678 0 sel[2]
<< properties >>
string FIXED_BBOX 0 0 10473 12617
<< end >>
