* NGSPICE file created from alu4bit.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

.subckt alu4bit A[0] A[1] A[2] A[3] B[0] B[1] B[2] B[3] VGND VPWR clk result[0] result[1]
+ result[2] result[3] rst sel[0] sel[1] sel[2]
XFILLER_0_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_062_ net12 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__buf_2
X_114_ _050_ _051_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ _050_ _051_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_112_ net7 _036_ _021_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_111_ net4 net8 VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__xnor2_1
X_110_ _035_ _040_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__o21ai_1
Xoutput13 net13 VGND VGND VPWR VPWR result[0] sky130_fd_sc_hd__buf_2
XFILLER_0_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR result[1] sky130_fd_sc_hd__clkbuf_4
X_099_ _037_ _038_ net3 VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__o21a_1
Xoutput15 net15 VGND VGND VPWR VPWR result[2] sky130_fd_sc_hd__clkbuf_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_098_ net7 _021_ _036_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__and3_1
Xoutput16 net16 VGND VGND VPWR VPWR result[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_097_ _021_ _036_ net7 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_096_ net5 net6 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_079_ _004_ _005_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__and2b_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_095_ _025_ _027_ _024_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__a21oi_2
X_078_ _005_ net10 _004_ net1 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nand4b_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_094_ _005_ net2 _004_ net10 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_077_ _018_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__clkbuf_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_093_ _015_ _019_ _032_ _033_ net9 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 A[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_076_ net9 _016_ _017_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ net2 net6 _015_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__a21oi_1
Xinput2 A[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_127_ clknet_1_1__leaf_clk _003_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
X_075_ net1 net5 _015_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a21o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 A[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_0_11_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_074_ _010_ _013_ _015_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__or3b_1
X_091_ _020_ _028_ _031_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__a21oi_1
X_126_ clknet_1_1__leaf_clk _002_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ _037_ _038_ net3 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 A[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_090_ net3 _011_ _012_ net2 _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_125_ clknet_1_0__leaf_clk _001_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_1
X_073_ _014_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__clkbuf_2
X_108_ _015_ _034_ _046_ _047_ net9 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 B[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_072_ _004_ net10 _005_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__or3_1
X_124_ clknet_1_0__leaf_clk _000_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_1
X_107_ net3 net7 _015_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 B[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_071_ net2 _011_ _012_ net1 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a22o_1
X_123_ _056_ _057_ _060_ _061_ net9 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__a311oi_1
X_106_ _020_ _042_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 B[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ _004_ net10 _005_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and3_1
XTAP_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 sel[0] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
X_122_ net4 net8 _015_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_105_ net4 _011_ _012_ net3 _044_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 B[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput11 sel[1] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
X_121_ net4 _012_ _058_ _059_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__a211oi_1
X_104_ net3 net7 _006_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__o22a_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 rst VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XTAP_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 sel[2] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
X_120_ net4 net8 _006_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_103_ net3 net7 _008_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_102_ _035_ _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ _039_ _040_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_100_ net3 _037_ _038_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_089_ net2 net6 _006_ _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__o22a_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_088_ net2 net6 _008_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ _026_ _027_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_086_ net1 net5 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ net10 _005_ _004_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ _024_ _025_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__or2b_1
XFILLER_0_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_068_ net1 net5 _006_ _009_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__o22a_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ _022_ _023_ net2 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_067_ net1 net5 _007_ _008_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a22oi_1
X_119_ _005_ net3 _004_ net10 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__and4b_1
XFILLER_0_6_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_083_ net2 _022_ _023_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__and3_1
X_118_ _004_ _050_ _005_ net10 VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_066_ net10 net11 net12 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__or3b_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_082_ net6 _021_ net5 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_065_ _004_ _005_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__or2b_1
X_117_ _049_ _052_ _053_ _055_ _007_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a311o_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_081_ net5 _021_ net6 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_064_ _004_ _005_ net10 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_116_ _035_ _040_ _054_ _048_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__o211a_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_080_ net12 net10 net11 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__nand3b_2
X_063_ net11 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__buf_2
X_115_ _052_ _053_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

