VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu4bit
  CLASS BLOCK ;
  FOREIGN alu4bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 52.365 BY 63.085 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 48.365 40.840 52.365 41.440 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 59.085 32.570 63.085 ;
    END
  END A[3]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 59.085 19.690 63.085 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 48.365 54.440 52.365 55.040 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END B[3]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.135 10.640 14.735 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.370 10.640 24.970 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.605 10.640 35.205 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.840 10.640 45.440 51.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.480 46.700 20.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 28.680 46.700 30.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 38.880 46.700 40.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 49.080 46.700 50.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.835 10.640 11.435 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.070 10.640 21.670 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.305 10.640 31.905 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.540 10.640 42.140 51.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.180 46.700 16.780 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 25.380 46.700 26.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 35.580 46.700 37.180 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 45.780 46.700 47.380 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END clk
  PIN result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 48.365 13.640 52.365 14.240 ;
    END
  END result[0]
  PIN result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END result[1]
  PIN result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END result[2]
  PIN result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 59.085 45.450 63.085 ;
    END
  END result[3]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END rst
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 59.085 6.810 63.085 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 48.365 27.240 52.365 27.840 ;
    END
  END sel[2]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 46.460 51.765 ;
      LAYER met1 ;
        RECT 0.070 10.640 51.910 51.920 ;
      LAYER met2 ;
        RECT 0.100 58.805 6.250 59.085 ;
        RECT 7.090 58.805 19.130 59.085 ;
        RECT 19.970 58.805 32.010 59.085 ;
        RECT 32.850 58.805 44.890 59.085 ;
        RECT 45.730 58.805 51.880 59.085 ;
        RECT 0.100 4.280 51.880 58.805 ;
        RECT 0.650 4.000 12.690 4.280 ;
        RECT 13.530 4.000 25.570 4.280 ;
        RECT 26.410 4.000 38.450 4.280 ;
        RECT 39.290 4.000 51.330 4.280 ;
      LAYER met3 ;
        RECT 4.400 54.040 47.965 54.905 ;
        RECT 4.000 41.840 48.365 54.040 ;
        RECT 4.400 40.440 47.965 41.840 ;
        RECT 4.000 28.240 48.365 40.440 ;
        RECT 4.400 26.840 47.965 28.240 ;
        RECT 4.000 14.640 48.365 26.840 ;
        RECT 4.400 13.240 47.965 14.640 ;
        RECT 4.000 10.715 48.365 13.240 ;
  END
END alu4bit
END LIBRARY

